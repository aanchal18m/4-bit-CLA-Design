magic
tech scmos
timestamp 1732025555
<< nwell >>
rect -21 -12 89 20
rect 96 -10 120 16
<< ntransistor >>
rect 107 -24 109 -19
rect -10 -30 -8 -25
rect 22 -35 24 -25
rect 33 -35 35 -25
rect 59 -35 61 -25
rect 70 -35 72 -25
<< ptransistor >>
rect -10 -6 -8 14
rect 0 -6 2 14
rect 22 -1 24 9
rect 59 -1 61 9
rect 107 0 109 10
<< ndiffusion >>
rect 106 -24 107 -19
rect 109 -24 110 -19
rect -11 -30 -10 -25
rect -8 -30 5 -25
rect 21 -35 22 -25
rect 24 -35 33 -25
rect 35 -35 40 -25
rect 57 -35 59 -25
rect 61 -35 70 -25
rect 72 -35 76 -25
<< pdiffusion >>
rect -11 -6 -10 14
rect -8 -6 0 14
rect 2 -6 5 14
rect 21 -1 22 9
rect 24 -1 40 9
rect 57 -1 59 9
rect 61 -1 76 9
rect 106 0 107 10
rect 109 0 110 10
<< ndcontact >>
rect 102 -24 106 -19
rect 110 -24 114 -19
rect -15 -30 -11 -25
rect 5 -30 9 -25
rect 17 -35 21 -25
rect 40 -35 44 -25
rect 53 -35 57 -25
rect 76 -35 80 -25
<< pdcontact >>
rect -15 -6 -11 14
rect 5 -6 9 14
rect 17 -1 21 9
rect 40 -1 44 9
rect 53 -1 57 9
rect 76 -1 80 9
rect 102 0 106 10
rect 110 0 114 10
<< polysilicon >>
rect -10 14 -8 17
rect 0 14 2 17
rect 22 9 24 13
rect 59 9 61 13
rect 107 10 109 14
rect -10 -25 -8 -6
rect 0 -22 2 -6
rect 22 -25 24 -1
rect 33 -25 35 -18
rect 59 -25 61 -1
rect 70 -25 72 -18
rect 107 -19 109 0
rect -10 -33 -8 -30
rect 107 -30 109 -24
rect 22 -38 24 -35
rect 33 -38 35 -35
rect 59 -38 61 -35
rect 70 -38 72 -35
<< polycontact >>
rect -14 -18 -10 -14
rect -4 -22 0 -18
rect 18 -18 22 -14
rect 55 -18 59 -14
rect 29 -22 33 -18
rect 103 -16 107 -12
rect 66 -22 70 -18
<< metal1 >>
rect -21 20 102 24
rect -15 14 -11 20
rect 17 9 21 20
rect 53 9 57 20
rect 95 16 120 20
rect 102 10 106 16
rect 5 -25 9 -6
rect 40 -14 44 -1
rect 76 -12 80 -1
rect 110 -12 114 0
rect 40 -18 55 -14
rect 76 -16 103 -12
rect 110 -16 122 -12
rect 40 -25 44 -18
rect 76 -25 80 -16
rect 110 -19 114 -16
rect -15 -41 -11 -30
rect 102 -33 106 -24
rect 17 -41 21 -35
rect 53 -41 57 -35
rect 98 -37 118 -33
rect 98 -41 102 -37
rect -15 -47 102 -41
<< labels >>
rlabel pdiffusion -5 4 -5 4 1 n1
rlabel pdcontact -13 4 -13 4 1 vdd
rlabel polycontact -12 -16 -12 -16 1 a
rlabel pdcontact 7 4 7 4 1 b
rlabel polycontact -2 -20 -2 -20 1 clk
rlabel ndcontact -13 -28 -13 -28 1 gnd
rlabel ndcontact 7 -28 7 -28 1 b
rlabel pdcontact 19 4 19 4 1 vdd
rlabel polycontact 31 -20 31 -20 1 b
rlabel ndcontact 19 -30 19 -30 1 gnd
rlabel ndiffusion 28 -30 28 -30 1 n2
rlabel ndcontact 42 -30 42 -30 1 c
rlabel pdcontact 42 4 42 4 1 c
rlabel ndcontact 78 -30 78 -30 1 n4
rlabel ndiffusion 65 -30 66 -30 1 n3
rlabel ndcontact 55 -30 55 -30 1 gnd
rlabel polycontact 68 -20 68 -20 1 clk
rlabel polycontact 57 -16 57 -16 1 c
rlabel pdcontact 55 3 55 3 1 vdd
rlabel pdcontact 78 4 78 4 1 n4
rlabel polycontact 20 -16 20 -16 1 clk
rlabel metal1 108 18 108 18 5 vdd
rlabel pdcontact 112 5 112 5 1 out
rlabel metal1 119 -14 119 -14 8 out
rlabel pdcontact 104 5 104 5 1 vdd
rlabel ndcontact 104 -22 104 -22 1 gnd
rlabel ndcontact 112 -22 112 -22 1 out
rlabel metal1 106 -35 106 -35 1 gnd
rlabel polycontact 105 -14 105 -14 1 n4
<< end >>
