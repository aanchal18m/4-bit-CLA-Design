magic
tech scmos
timestamp 1732053798
<< nwell >>
rect -1129 803 -1077 806
rect -1188 776 -1164 802
rect -1155 777 -1077 803
rect -1043 787 -991 806
rect -955 789 -920 797
rect -1129 771 -1077 777
rect -1071 771 -991 787
rect -1071 761 -1047 771
rect -985 761 -961 787
rect -955 764 -893 789
rect -917 763 -893 764
rect -997 683 -945 718
rect -939 673 -915 699
rect -654 613 -602 648
rect -596 603 -572 629
rect -1131 591 -1079 594
rect -1190 564 -1166 590
rect -1157 565 -1079 591
rect -1045 575 -993 594
rect -957 577 -922 585
rect -1131 559 -1079 565
rect -1073 559 -993 575
rect -1073 549 -1049 559
rect -987 549 -963 575
rect -957 552 -895 577
rect -919 551 -895 552
rect -658 527 -596 547
rect -523 543 -462 563
rect -658 523 -571 527
rect -658 512 -568 523
rect -999 471 -947 506
rect -592 497 -568 512
rect -523 517 -433 543
rect -523 511 -462 517
rect -941 461 -917 487
rect -661 405 -596 425
rect -241 405 -189 408
rect -661 401 -574 405
rect -661 390 -571 401
rect -1132 376 -1080 379
rect -1191 349 -1167 375
rect -1158 350 -1080 376
rect -1046 360 -994 379
rect -595 375 -571 390
rect -300 378 -276 404
rect -267 379 -189 405
rect -155 389 -103 408
rect -67 391 -32 399
rect -241 373 -189 379
rect -183 373 -103 389
rect -958 362 -923 370
rect -183 363 -159 373
rect -97 363 -73 389
rect -67 366 -5 391
rect -29 365 -5 366
rect -1132 344 -1080 350
rect -1074 344 -994 360
rect -1074 334 -1050 344
rect -988 334 -964 360
rect -958 337 -896 362
rect -920 336 -896 337
rect -1000 256 -948 291
rect -942 246 -918 272
rect -672 256 -620 291
rect -241 288 -189 291
rect -614 246 -590 272
rect -562 249 -501 262
rect -300 261 -276 287
rect -267 262 -189 288
rect -155 272 -103 291
rect -67 274 -32 282
rect -241 256 -189 262
rect -183 256 -103 272
rect -562 223 -472 249
rect -183 246 -159 256
rect -97 246 -73 272
rect -67 249 -5 274
rect -29 248 -5 249
rect -562 217 -501 223
rect -676 170 -614 190
rect -676 166 -589 170
rect -243 168 -191 171
rect -676 155 -586 166
rect -1129 148 -1077 151
rect -1188 121 -1164 147
rect -1155 122 -1077 148
rect -1043 132 -991 151
rect -955 134 -920 142
rect -610 140 -586 155
rect -302 141 -278 167
rect -269 142 -191 168
rect -157 152 -105 171
rect -69 154 -34 162
rect -243 136 -191 142
rect -185 136 -105 152
rect -1129 116 -1077 122
rect -1071 116 -991 132
rect -1071 106 -1047 116
rect -985 106 -961 132
rect -955 109 -893 134
rect -185 126 -161 136
rect -99 126 -75 152
rect -69 129 -7 154
rect -31 128 -7 129
rect -917 108 -893 109
rect -997 28 -945 63
rect -939 18 -915 44
rect -675 35 -623 70
rect -580 58 -545 66
rect -617 25 -593 51
rect -580 33 -518 58
rect -243 51 -191 54
rect -542 32 -518 33
rect -302 24 -278 50
rect -269 25 -191 51
rect -157 35 -105 54
rect -69 37 -34 45
rect -243 19 -191 25
rect -185 19 -105 35
rect -185 9 -161 19
rect -99 9 -75 35
rect -69 12 -7 37
rect -31 11 -7 12
<< ntransistor >>
rect -1177 762 -1175 767
rect -1144 763 -1142 768
rect -1113 741 -1110 751
rect -1099 741 -1096 751
rect -1060 747 -1058 752
rect -1027 741 -1024 751
rect -1013 741 -1010 751
rect -974 747 -972 752
rect -906 749 -904 754
rect -944 742 -942 747
rect -933 742 -931 747
rect -981 653 -978 663
rect -967 653 -964 663
rect -928 659 -926 664
rect -638 583 -635 593
rect -624 583 -621 593
rect -585 589 -583 594
rect -1179 550 -1177 555
rect -1146 551 -1144 556
rect -1115 529 -1112 539
rect -1101 529 -1098 539
rect -1062 535 -1060 540
rect -1029 529 -1026 539
rect -1015 529 -1012 539
rect -976 535 -974 540
rect -908 537 -906 542
rect -946 530 -944 535
rect -935 530 -933 535
rect -642 469 -639 484
rect -628 469 -625 484
rect -613 469 -610 484
rect -581 483 -579 488
rect -446 503 -444 508
rect -512 477 -510 482
rect -501 477 -499 482
rect -490 477 -488 482
rect -480 477 -478 482
rect -983 441 -980 451
rect -969 441 -966 451
rect -930 447 -928 452
rect -1180 335 -1178 340
rect -1147 336 -1145 341
rect -1116 314 -1113 324
rect -1102 314 -1099 324
rect -1063 320 -1061 325
rect -1030 314 -1027 324
rect -1016 314 -1013 324
rect -977 320 -975 325
rect -645 342 -642 362
rect -631 342 -628 362
rect -620 342 -617 362
rect -611 342 -608 362
rect -584 361 -582 366
rect -289 364 -287 369
rect -256 365 -254 370
rect -225 343 -222 353
rect -211 343 -208 353
rect -172 349 -170 354
rect -139 343 -136 353
rect -125 343 -122 353
rect -86 349 -84 354
rect -18 351 -16 356
rect -56 344 -54 349
rect -45 344 -43 349
rect -909 322 -907 327
rect -947 315 -945 320
rect -936 315 -934 320
rect -984 226 -981 236
rect -970 226 -967 236
rect -931 232 -929 237
rect -656 226 -653 236
rect -642 226 -639 236
rect -603 232 -601 237
rect -289 247 -287 252
rect -256 248 -254 253
rect -225 226 -222 236
rect -211 226 -208 236
rect -172 232 -170 237
rect -139 226 -136 236
rect -125 226 -122 236
rect -86 232 -84 237
rect -18 234 -16 239
rect -56 227 -54 232
rect -45 227 -43 232
rect -485 209 -483 214
rect -551 185 -549 189
rect -540 185 -538 189
rect -527 185 -525 189
rect -1177 107 -1175 112
rect -1144 108 -1142 113
rect -1113 86 -1110 96
rect -1099 86 -1096 96
rect -1060 92 -1058 97
rect -1027 86 -1024 96
rect -1013 86 -1010 96
rect -974 92 -972 97
rect -660 112 -657 127
rect -646 112 -643 127
rect -631 112 -628 127
rect -599 126 -597 131
rect -291 127 -289 132
rect -258 128 -256 133
rect -227 106 -224 116
rect -213 106 -210 116
rect -174 112 -172 117
rect -141 106 -138 116
rect -127 106 -124 116
rect -88 112 -86 117
rect -20 114 -18 119
rect -58 107 -56 112
rect -47 107 -45 112
rect -906 94 -904 99
rect -944 87 -942 92
rect -933 87 -931 92
rect -531 18 -529 23
rect -981 -2 -978 8
rect -967 -2 -964 8
rect -928 4 -926 9
rect -659 5 -656 15
rect -645 5 -642 15
rect -606 11 -604 16
rect -569 11 -567 16
rect -558 11 -556 16
rect -291 10 -289 15
rect -258 11 -256 16
rect -227 -11 -224 -1
rect -213 -11 -210 -1
rect -174 -5 -172 0
rect -141 -11 -138 -1
rect -127 -11 -124 -1
rect -88 -5 -86 0
rect -20 -3 -18 2
rect -58 -10 -56 -5
rect -47 -10 -45 -5
<< ptransistor >>
rect -1177 786 -1175 796
rect -1144 787 -1142 797
rect -1113 788 -1110 798
rect -1099 788 -1096 798
rect -1027 788 -1024 798
rect -1013 788 -1010 798
rect -1060 771 -1058 781
rect -974 771 -972 781
rect -944 771 -942 791
rect -933 771 -931 791
rect -906 773 -904 783
rect -981 700 -978 710
rect -967 700 -964 710
rect -928 683 -926 693
rect -638 630 -635 640
rect -624 630 -621 640
rect -585 613 -583 623
rect -1179 574 -1177 584
rect -1146 575 -1144 585
rect -1115 576 -1112 586
rect -1101 576 -1098 586
rect -1029 576 -1026 586
rect -1015 576 -1012 586
rect -1062 559 -1060 569
rect -976 559 -974 569
rect -946 559 -944 579
rect -935 559 -933 579
rect -908 561 -906 571
rect -642 529 -639 539
rect -628 529 -625 539
rect -613 529 -610 539
rect -983 488 -980 498
rect -969 488 -966 498
rect -512 517 -510 557
rect -501 517 -499 557
rect -490 517 -488 557
rect -480 517 -478 557
rect -446 527 -444 537
rect -581 507 -579 517
rect -930 471 -928 481
rect -645 407 -642 417
rect -631 407 -628 417
rect -620 407 -617 417
rect -611 407 -608 417
rect -1180 359 -1178 369
rect -1147 360 -1145 370
rect -1116 361 -1113 371
rect -1102 361 -1099 371
rect -1030 361 -1027 371
rect -1016 361 -1013 371
rect -1063 344 -1061 354
rect -977 344 -975 354
rect -947 344 -945 364
rect -936 344 -934 364
rect -584 385 -582 395
rect -289 388 -287 398
rect -256 389 -254 399
rect -225 390 -222 400
rect -211 390 -208 400
rect -139 390 -136 400
rect -125 390 -122 400
rect -909 346 -907 356
rect -172 373 -170 383
rect -86 373 -84 383
rect -56 373 -54 393
rect -45 373 -43 393
rect -18 375 -16 385
rect -984 273 -981 283
rect -970 273 -967 283
rect -656 273 -653 283
rect -642 273 -639 283
rect -931 256 -929 266
rect -289 271 -287 281
rect -256 272 -254 282
rect -225 273 -222 283
rect -211 273 -208 283
rect -139 273 -136 283
rect -125 273 -122 283
rect -603 256 -601 266
rect -551 224 -549 254
rect -540 224 -538 254
rect -527 224 -525 254
rect -485 233 -483 243
rect -172 256 -170 266
rect -86 256 -84 266
rect -56 256 -54 276
rect -45 256 -43 276
rect -18 258 -16 268
rect -660 172 -657 182
rect -646 172 -643 182
rect -631 172 -628 182
rect -1177 131 -1175 141
rect -1144 132 -1142 142
rect -1113 133 -1110 143
rect -1099 133 -1096 143
rect -1027 133 -1024 143
rect -1013 133 -1010 143
rect -1060 116 -1058 126
rect -974 116 -972 126
rect -944 116 -942 136
rect -933 116 -931 136
rect -906 118 -904 128
rect -599 150 -597 160
rect -291 151 -289 161
rect -258 152 -256 162
rect -227 153 -224 163
rect -213 153 -210 163
rect -141 153 -138 163
rect -127 153 -124 163
rect -174 136 -172 146
rect -88 136 -86 146
rect -58 136 -56 156
rect -47 136 -45 156
rect -20 138 -18 148
rect -981 45 -978 55
rect -967 45 -964 55
rect -659 52 -656 62
rect -645 52 -642 62
rect -928 28 -926 38
rect -606 35 -604 45
rect -569 40 -567 60
rect -558 40 -556 60
rect -531 42 -529 52
rect -291 34 -289 44
rect -258 35 -256 45
rect -227 36 -224 46
rect -213 36 -210 46
rect -141 36 -138 46
rect -127 36 -124 46
rect -174 19 -172 29
rect -88 19 -86 29
rect -58 19 -56 39
rect -47 19 -45 39
rect -20 21 -18 31
<< ndiffusion >>
rect -1178 762 -1177 767
rect -1175 762 -1174 767
rect -1145 763 -1144 768
rect -1142 763 -1141 768
rect -1116 741 -1113 751
rect -1110 741 -1099 751
rect -1096 741 -1090 751
rect -1061 747 -1060 752
rect -1058 747 -1057 752
rect -1030 741 -1027 751
rect -1024 741 -1013 751
rect -1010 741 -1004 751
rect -975 747 -974 752
rect -972 747 -971 752
rect -907 749 -906 754
rect -904 749 -903 754
rect -945 742 -944 747
rect -942 742 -940 747
rect -936 742 -933 747
rect -931 742 -930 747
rect -984 653 -981 663
rect -978 653 -967 663
rect -964 653 -958 663
rect -929 659 -928 664
rect -926 659 -925 664
rect -641 583 -638 593
rect -635 583 -624 593
rect -621 583 -615 593
rect -586 589 -585 594
rect -583 589 -582 594
rect -1180 550 -1179 555
rect -1177 550 -1176 555
rect -1147 551 -1146 556
rect -1144 551 -1143 556
rect -1118 529 -1115 539
rect -1112 529 -1101 539
rect -1098 529 -1092 539
rect -1063 535 -1062 540
rect -1060 535 -1059 540
rect -1032 529 -1029 539
rect -1026 529 -1015 539
rect -1012 529 -1006 539
rect -977 535 -976 540
rect -974 535 -973 540
rect -909 537 -908 542
rect -906 537 -905 542
rect -947 530 -946 535
rect -944 530 -942 535
rect -938 530 -935 535
rect -933 530 -932 535
rect -646 469 -642 484
rect -639 469 -628 484
rect -625 469 -613 484
rect -610 469 -607 484
rect -582 483 -581 488
rect -579 483 -578 488
rect -447 503 -446 508
rect -444 503 -443 508
rect -513 477 -512 482
rect -510 477 -507 482
rect -503 477 -501 482
rect -499 477 -495 482
rect -491 477 -490 482
rect -488 477 -486 482
rect -482 477 -480 482
rect -478 477 -477 482
rect -986 441 -983 451
rect -980 441 -969 451
rect -966 441 -960 451
rect -931 447 -930 452
rect -928 447 -927 452
rect -1181 335 -1180 340
rect -1178 335 -1177 340
rect -1148 336 -1147 341
rect -1145 336 -1144 341
rect -1119 314 -1116 324
rect -1113 314 -1102 324
rect -1099 314 -1093 324
rect -1064 320 -1063 325
rect -1061 320 -1060 325
rect -1033 314 -1030 324
rect -1027 314 -1016 324
rect -1013 314 -1007 324
rect -978 320 -977 325
rect -975 320 -974 325
rect -649 342 -645 362
rect -642 342 -631 362
rect -628 342 -620 362
rect -617 342 -611 362
rect -608 342 -605 362
rect -585 361 -584 366
rect -582 361 -581 366
rect -290 364 -289 369
rect -287 364 -286 369
rect -257 365 -256 370
rect -254 365 -253 370
rect -228 343 -225 353
rect -222 343 -211 353
rect -208 343 -202 353
rect -173 349 -172 354
rect -170 349 -169 354
rect -142 343 -139 353
rect -136 343 -125 353
rect -122 343 -116 353
rect -87 349 -86 354
rect -84 349 -83 354
rect -19 351 -18 356
rect -16 351 -15 356
rect -57 344 -56 349
rect -54 344 -52 349
rect -48 344 -45 349
rect -43 344 -42 349
rect -910 322 -909 327
rect -907 322 -906 327
rect -948 315 -947 320
rect -945 315 -943 320
rect -939 315 -936 320
rect -934 315 -933 320
rect -987 226 -984 236
rect -981 226 -970 236
rect -967 226 -961 236
rect -932 232 -931 237
rect -929 232 -928 237
rect -659 226 -656 236
rect -653 226 -642 236
rect -639 226 -633 236
rect -604 232 -603 237
rect -601 232 -600 237
rect -290 247 -289 252
rect -287 247 -286 252
rect -257 248 -256 253
rect -254 248 -253 253
rect -228 226 -225 236
rect -222 226 -211 236
rect -208 226 -202 236
rect -173 232 -172 237
rect -170 232 -169 237
rect -142 226 -139 236
rect -136 226 -125 236
rect -122 226 -116 236
rect -87 232 -86 237
rect -84 232 -83 237
rect -19 234 -18 239
rect -16 234 -15 239
rect -57 227 -56 232
rect -54 227 -52 232
rect -48 227 -45 232
rect -43 227 -42 232
rect -486 209 -485 214
rect -483 209 -482 214
rect -552 185 -551 189
rect -549 185 -546 189
rect -542 185 -540 189
rect -538 185 -534 189
rect -530 185 -527 189
rect -525 185 -516 189
rect -1178 107 -1177 112
rect -1175 107 -1174 112
rect -1145 108 -1144 113
rect -1142 108 -1141 113
rect -1116 86 -1113 96
rect -1110 86 -1099 96
rect -1096 86 -1090 96
rect -1061 92 -1060 97
rect -1058 92 -1057 97
rect -1030 86 -1027 96
rect -1024 86 -1013 96
rect -1010 86 -1004 96
rect -975 92 -974 97
rect -972 92 -971 97
rect -664 112 -660 127
rect -657 112 -646 127
rect -643 112 -631 127
rect -628 112 -625 127
rect -600 126 -599 131
rect -597 126 -596 131
rect -292 127 -291 132
rect -289 127 -288 132
rect -259 128 -258 133
rect -256 128 -255 133
rect -230 106 -227 116
rect -224 106 -213 116
rect -210 106 -204 116
rect -175 112 -174 117
rect -172 112 -171 117
rect -144 106 -141 116
rect -138 106 -127 116
rect -124 106 -118 116
rect -89 112 -88 117
rect -86 112 -85 117
rect -21 114 -20 119
rect -18 114 -17 119
rect -59 107 -58 112
rect -56 107 -54 112
rect -50 107 -47 112
rect -45 107 -44 112
rect -907 94 -906 99
rect -904 94 -903 99
rect -945 87 -944 92
rect -942 87 -940 92
rect -936 87 -933 92
rect -931 87 -930 92
rect -532 18 -531 23
rect -529 18 -528 23
rect -984 -2 -981 8
rect -978 -2 -967 8
rect -964 -2 -958 8
rect -929 4 -928 9
rect -926 4 -925 9
rect -662 5 -659 15
rect -656 5 -645 15
rect -642 5 -636 15
rect -607 11 -606 16
rect -604 11 -603 16
rect -570 11 -569 16
rect -567 11 -565 16
rect -561 11 -558 16
rect -556 11 -555 16
rect -292 10 -291 15
rect -289 10 -288 15
rect -259 11 -258 16
rect -256 11 -255 16
rect -230 -11 -227 -1
rect -224 -11 -213 -1
rect -210 -11 -204 -1
rect -175 -5 -174 0
rect -172 -5 -171 0
rect -144 -11 -141 -1
rect -138 -11 -127 -1
rect -124 -11 -118 -1
rect -89 -5 -88 0
rect -86 -5 -85 0
rect -21 -3 -20 2
rect -18 -3 -17 2
rect -59 -10 -58 -5
rect -56 -10 -54 -5
rect -50 -10 -47 -5
rect -45 -10 -44 -5
<< pdiffusion >>
rect -1178 786 -1177 796
rect -1175 786 -1174 796
rect -1145 787 -1144 797
rect -1142 787 -1141 797
rect -1116 788 -1113 798
rect -1110 788 -1107 798
rect -1102 788 -1099 798
rect -1096 788 -1090 798
rect -1030 788 -1027 798
rect -1024 788 -1021 798
rect -1016 788 -1013 798
rect -1010 788 -1004 798
rect -1061 771 -1060 781
rect -1058 771 -1057 781
rect -975 771 -974 781
rect -972 771 -971 781
rect -945 771 -944 791
rect -942 771 -933 791
rect -931 771 -930 791
rect -907 773 -906 783
rect -904 773 -903 783
rect -984 700 -981 710
rect -978 700 -975 710
rect -970 700 -967 710
rect -964 700 -958 710
rect -929 683 -928 693
rect -926 683 -925 693
rect -641 630 -638 640
rect -635 630 -632 640
rect -627 630 -624 640
rect -621 630 -615 640
rect -586 613 -585 623
rect -583 613 -582 623
rect -1180 574 -1179 584
rect -1177 574 -1176 584
rect -1147 575 -1146 585
rect -1144 575 -1143 585
rect -1118 576 -1115 586
rect -1112 576 -1109 586
rect -1104 576 -1101 586
rect -1098 576 -1092 586
rect -1032 576 -1029 586
rect -1026 576 -1023 586
rect -1018 576 -1015 586
rect -1012 576 -1006 586
rect -1063 559 -1062 569
rect -1060 559 -1059 569
rect -977 559 -976 569
rect -974 559 -973 569
rect -947 559 -946 579
rect -944 559 -935 579
rect -933 559 -932 579
rect -909 561 -908 571
rect -906 561 -905 571
rect -645 529 -642 539
rect -639 529 -636 539
rect -631 529 -628 539
rect -625 529 -619 539
rect -614 529 -613 539
rect -610 529 -607 539
rect -986 488 -983 498
rect -980 488 -977 498
rect -972 488 -969 498
rect -966 488 -960 498
rect -513 517 -512 557
rect -510 517 -501 557
rect -499 517 -490 557
rect -488 517 -480 557
rect -478 517 -477 557
rect -447 527 -446 537
rect -444 527 -443 537
rect -582 507 -581 517
rect -579 507 -578 517
rect -931 471 -930 481
rect -928 471 -927 481
rect -648 407 -645 417
rect -642 407 -639 417
rect -634 407 -631 417
rect -628 407 -626 417
rect -622 407 -620 417
rect -617 407 -616 417
rect -612 407 -611 417
rect -608 407 -606 417
rect -1181 359 -1180 369
rect -1178 359 -1177 369
rect -1148 360 -1147 370
rect -1145 360 -1144 370
rect -1119 361 -1116 371
rect -1113 361 -1110 371
rect -1105 361 -1102 371
rect -1099 361 -1093 371
rect -1033 361 -1030 371
rect -1027 361 -1024 371
rect -1019 361 -1016 371
rect -1013 361 -1007 371
rect -1064 344 -1063 354
rect -1061 344 -1060 354
rect -978 344 -977 354
rect -975 344 -974 354
rect -948 344 -947 364
rect -945 344 -936 364
rect -934 344 -933 364
rect -585 385 -584 395
rect -582 385 -581 395
rect -290 388 -289 398
rect -287 388 -286 398
rect -257 389 -256 399
rect -254 389 -253 399
rect -228 390 -225 400
rect -222 390 -219 400
rect -214 390 -211 400
rect -208 390 -202 400
rect -142 390 -139 400
rect -136 390 -133 400
rect -128 390 -125 400
rect -122 390 -116 400
rect -910 346 -909 356
rect -907 346 -906 356
rect -173 373 -172 383
rect -170 373 -169 383
rect -87 373 -86 383
rect -84 373 -83 383
rect -57 373 -56 393
rect -54 373 -45 393
rect -43 373 -42 393
rect -19 375 -18 385
rect -16 375 -15 385
rect -987 273 -984 283
rect -981 273 -978 283
rect -973 273 -970 283
rect -967 273 -961 283
rect -659 273 -656 283
rect -653 273 -650 283
rect -645 273 -642 283
rect -639 273 -633 283
rect -932 256 -931 266
rect -929 256 -928 266
rect -290 271 -289 281
rect -287 271 -286 281
rect -257 272 -256 282
rect -254 272 -253 282
rect -228 273 -225 283
rect -222 273 -219 283
rect -214 273 -211 283
rect -208 273 -202 283
rect -142 273 -139 283
rect -136 273 -133 283
rect -128 273 -125 283
rect -122 273 -116 283
rect -604 256 -603 266
rect -601 256 -600 266
rect -552 224 -551 254
rect -549 224 -540 254
rect -538 224 -527 254
rect -525 224 -516 254
rect -486 233 -485 243
rect -483 233 -482 243
rect -173 256 -172 266
rect -170 256 -169 266
rect -87 256 -86 266
rect -84 256 -83 266
rect -57 256 -56 276
rect -54 256 -45 276
rect -43 256 -42 276
rect -19 258 -18 268
rect -16 258 -15 268
rect -663 172 -660 182
rect -657 172 -654 182
rect -649 172 -646 182
rect -643 172 -637 182
rect -632 172 -631 182
rect -628 172 -625 182
rect -1178 131 -1177 141
rect -1175 131 -1174 141
rect -1145 132 -1144 142
rect -1142 132 -1141 142
rect -1116 133 -1113 143
rect -1110 133 -1107 143
rect -1102 133 -1099 143
rect -1096 133 -1090 143
rect -1030 133 -1027 143
rect -1024 133 -1021 143
rect -1016 133 -1013 143
rect -1010 133 -1004 143
rect -1061 116 -1060 126
rect -1058 116 -1057 126
rect -975 116 -974 126
rect -972 116 -971 126
rect -945 116 -944 136
rect -942 116 -933 136
rect -931 116 -930 136
rect -907 118 -906 128
rect -904 118 -903 128
rect -600 150 -599 160
rect -597 150 -596 160
rect -292 151 -291 161
rect -289 151 -288 161
rect -259 152 -258 162
rect -256 152 -255 162
rect -230 153 -227 163
rect -224 153 -221 163
rect -216 153 -213 163
rect -210 153 -204 163
rect -144 153 -141 163
rect -138 153 -135 163
rect -130 153 -127 163
rect -124 153 -118 163
rect -175 136 -174 146
rect -172 136 -171 146
rect -89 136 -88 146
rect -86 136 -85 146
rect -59 136 -58 156
rect -56 136 -47 156
rect -45 136 -44 156
rect -21 138 -20 148
rect -18 138 -17 148
rect -984 45 -981 55
rect -978 45 -975 55
rect -970 45 -967 55
rect -964 45 -958 55
rect -662 52 -659 62
rect -656 52 -653 62
rect -648 52 -645 62
rect -642 52 -636 62
rect -929 28 -928 38
rect -926 28 -925 38
rect -607 35 -606 45
rect -604 35 -603 45
rect -570 40 -569 60
rect -567 40 -558 60
rect -556 40 -555 60
rect -532 42 -531 52
rect -529 42 -528 52
rect -292 34 -291 44
rect -289 34 -288 44
rect -259 35 -258 45
rect -256 35 -255 45
rect -230 36 -227 46
rect -224 36 -221 46
rect -216 36 -213 46
rect -210 36 -204 46
rect -144 36 -141 46
rect -138 36 -135 46
rect -130 36 -127 46
rect -124 36 -118 46
rect -175 19 -174 29
rect -172 19 -171 29
rect -89 19 -88 29
rect -86 19 -85 29
rect -59 19 -58 39
rect -56 19 -47 39
rect -45 19 -44 39
rect -21 21 -20 31
rect -18 21 -17 31
<< ndcontact >>
rect -1182 762 -1178 767
rect -1174 762 -1170 767
rect -1149 763 -1145 768
rect -1141 763 -1137 768
rect -1121 741 -1116 751
rect -1090 741 -1085 751
rect -1065 747 -1061 752
rect -1057 747 -1053 752
rect -1035 741 -1030 751
rect -1004 741 -999 751
rect -979 747 -975 752
rect -971 747 -967 752
rect -911 749 -907 754
rect -903 749 -899 754
rect -949 742 -945 747
rect -940 742 -936 747
rect -930 742 -926 747
rect -989 653 -984 663
rect -958 653 -953 663
rect -933 659 -929 664
rect -925 659 -921 664
rect -646 583 -641 593
rect -615 583 -610 593
rect -590 589 -586 594
rect -582 589 -578 594
rect -1184 550 -1180 555
rect -1176 550 -1172 555
rect -1151 551 -1147 556
rect -1143 551 -1139 556
rect -1123 529 -1118 539
rect -1092 529 -1087 539
rect -1067 535 -1063 540
rect -1059 535 -1055 540
rect -1037 529 -1032 539
rect -1006 529 -1001 539
rect -981 535 -977 540
rect -973 535 -969 540
rect -913 537 -909 542
rect -905 537 -901 542
rect -951 530 -947 535
rect -942 530 -938 535
rect -932 530 -928 535
rect -650 469 -646 484
rect -607 469 -603 484
rect -586 483 -582 488
rect -578 483 -574 488
rect -451 503 -447 508
rect -443 503 -439 508
rect -517 477 -513 482
rect -507 477 -503 482
rect -495 477 -491 482
rect -486 477 -482 482
rect -477 477 -471 482
rect -991 441 -986 451
rect -960 441 -955 451
rect -935 447 -931 452
rect -927 447 -923 452
rect -1185 335 -1181 340
rect -1177 335 -1173 340
rect -1152 336 -1148 341
rect -1144 336 -1140 341
rect -1124 314 -1119 324
rect -1093 314 -1088 324
rect -1068 320 -1064 325
rect -1060 320 -1056 325
rect -1038 314 -1033 324
rect -1007 314 -1002 324
rect -982 320 -978 325
rect -974 320 -970 325
rect -653 342 -649 362
rect -605 342 -601 362
rect -589 361 -585 366
rect -581 361 -577 366
rect -294 364 -290 369
rect -286 364 -282 369
rect -261 365 -257 370
rect -253 365 -249 370
rect -233 343 -228 353
rect -202 343 -197 353
rect -177 349 -173 354
rect -169 349 -165 354
rect -147 343 -142 353
rect -116 343 -111 353
rect -91 349 -87 354
rect -83 349 -79 354
rect -23 351 -19 356
rect -15 351 -11 356
rect -61 344 -57 349
rect -52 344 -48 349
rect -42 344 -38 349
rect -914 322 -910 327
rect -906 322 -902 327
rect -952 315 -948 320
rect -943 315 -939 320
rect -933 315 -929 320
rect -992 226 -987 236
rect -961 226 -956 236
rect -936 232 -932 237
rect -928 232 -924 237
rect -664 226 -659 236
rect -633 226 -628 236
rect -608 232 -604 237
rect -600 232 -596 237
rect -294 247 -290 252
rect -286 247 -282 252
rect -261 248 -257 253
rect -253 248 -249 253
rect -233 226 -228 236
rect -202 226 -197 236
rect -177 232 -173 237
rect -169 232 -165 237
rect -147 226 -142 236
rect -116 226 -111 236
rect -91 232 -87 237
rect -83 232 -79 237
rect -23 234 -19 239
rect -15 234 -11 239
rect -61 227 -57 232
rect -52 227 -48 232
rect -42 227 -38 232
rect -490 209 -486 214
rect -482 209 -478 214
rect -556 185 -552 189
rect -546 185 -542 189
rect -534 185 -530 189
rect -516 185 -510 189
rect -1182 107 -1178 112
rect -1174 107 -1170 112
rect -1149 108 -1145 113
rect -1141 108 -1137 113
rect -1121 86 -1116 96
rect -1090 86 -1085 96
rect -1065 92 -1061 97
rect -1057 92 -1053 97
rect -1035 86 -1030 96
rect -1004 86 -999 96
rect -979 92 -975 97
rect -971 92 -967 97
rect -668 112 -664 127
rect -625 112 -621 127
rect -604 126 -600 131
rect -596 126 -592 131
rect -296 127 -292 132
rect -288 127 -284 132
rect -263 128 -259 133
rect -255 128 -251 133
rect -235 106 -230 116
rect -204 106 -199 116
rect -179 112 -175 117
rect -171 112 -167 117
rect -149 106 -144 116
rect -118 106 -113 116
rect -93 112 -89 117
rect -85 112 -81 117
rect -25 114 -21 119
rect -17 114 -13 119
rect -63 107 -59 112
rect -54 107 -50 112
rect -44 107 -40 112
rect -911 94 -907 99
rect -903 94 -899 99
rect -949 87 -945 92
rect -940 87 -936 92
rect -930 87 -926 92
rect -536 18 -532 23
rect -528 18 -524 23
rect -989 -2 -984 8
rect -958 -2 -953 8
rect -933 4 -929 9
rect -925 4 -921 9
rect -667 5 -662 15
rect -636 5 -631 15
rect -611 11 -607 16
rect -603 11 -599 16
rect -574 11 -570 16
rect -565 11 -561 16
rect -555 11 -551 16
rect -296 10 -292 15
rect -288 10 -284 15
rect -263 11 -259 16
rect -255 11 -251 16
rect -235 -11 -230 -1
rect -204 -11 -199 -1
rect -179 -5 -175 0
rect -171 -5 -167 0
rect -149 -11 -144 -1
rect -118 -11 -113 -1
rect -93 -5 -89 0
rect -85 -5 -81 0
rect -25 -3 -21 2
rect -17 -3 -13 2
rect -63 -10 -59 -5
rect -54 -10 -50 -5
rect -44 -10 -40 -5
<< pdcontact >>
rect -1182 786 -1178 796
rect -1174 786 -1170 796
rect -1149 787 -1145 797
rect -1141 787 -1137 797
rect -1121 788 -1116 798
rect -1107 788 -1102 798
rect -1090 788 -1085 798
rect -1035 788 -1030 798
rect -1021 788 -1016 798
rect -1004 788 -999 798
rect -1065 771 -1061 781
rect -1057 771 -1053 781
rect -979 771 -975 781
rect -971 771 -967 781
rect -949 771 -945 791
rect -930 771 -926 791
rect -911 773 -907 783
rect -903 773 -899 783
rect -989 700 -984 710
rect -975 700 -970 710
rect -958 700 -953 710
rect -933 683 -929 693
rect -925 683 -921 693
rect -646 630 -641 640
rect -632 630 -627 640
rect -615 630 -610 640
rect -590 613 -586 623
rect -582 613 -578 623
rect -1184 574 -1180 584
rect -1176 574 -1172 584
rect -1151 575 -1147 585
rect -1143 575 -1139 585
rect -1123 576 -1118 586
rect -1109 576 -1104 586
rect -1092 576 -1087 586
rect -1037 576 -1032 586
rect -1023 576 -1018 586
rect -1006 576 -1001 586
rect -1067 559 -1063 569
rect -1059 559 -1055 569
rect -981 559 -977 569
rect -973 559 -969 569
rect -951 559 -947 579
rect -932 559 -928 579
rect -913 561 -909 571
rect -905 561 -901 571
rect -650 529 -645 539
rect -636 529 -631 539
rect -619 529 -614 539
rect -607 529 -603 539
rect -991 488 -986 498
rect -977 488 -972 498
rect -960 488 -955 498
rect -517 517 -513 557
rect -477 517 -471 557
rect -451 527 -447 537
rect -443 527 -439 537
rect -586 507 -582 517
rect -578 507 -574 517
rect -935 471 -931 481
rect -927 471 -923 481
rect -653 407 -648 417
rect -639 407 -634 417
rect -626 407 -622 417
rect -616 407 -612 417
rect -606 407 -602 417
rect -1185 359 -1181 369
rect -1177 359 -1173 369
rect -1152 360 -1148 370
rect -1144 360 -1140 370
rect -1124 361 -1119 371
rect -1110 361 -1105 371
rect -1093 361 -1088 371
rect -1038 361 -1033 371
rect -1024 361 -1019 371
rect -1007 361 -1002 371
rect -1068 344 -1064 354
rect -1060 344 -1056 354
rect -982 344 -978 354
rect -974 344 -970 354
rect -952 344 -948 364
rect -933 344 -929 364
rect -589 385 -585 395
rect -581 385 -577 395
rect -294 388 -290 398
rect -286 388 -282 398
rect -261 389 -257 399
rect -253 389 -249 399
rect -233 390 -228 400
rect -219 390 -214 400
rect -202 390 -197 400
rect -147 390 -142 400
rect -133 390 -128 400
rect -116 390 -111 400
rect -914 346 -910 356
rect -906 346 -902 356
rect -177 373 -173 383
rect -169 373 -165 383
rect -91 373 -87 383
rect -83 373 -79 383
rect -61 373 -57 393
rect -42 373 -38 393
rect -23 375 -19 385
rect -15 375 -11 385
rect -992 273 -987 283
rect -978 273 -973 283
rect -961 273 -956 283
rect -664 273 -659 283
rect -650 273 -645 283
rect -633 273 -628 283
rect -936 256 -932 266
rect -928 256 -924 266
rect -294 271 -290 281
rect -286 271 -282 281
rect -261 272 -257 282
rect -253 272 -249 282
rect -233 273 -228 283
rect -219 273 -214 283
rect -202 273 -197 283
rect -147 273 -142 283
rect -133 273 -128 283
rect -116 273 -111 283
rect -608 256 -604 266
rect -600 256 -596 266
rect -556 224 -552 254
rect -516 224 -510 254
rect -490 233 -486 243
rect -482 233 -478 243
rect -177 256 -173 266
rect -169 256 -165 266
rect -91 256 -87 266
rect -83 256 -79 266
rect -61 256 -57 276
rect -42 256 -38 276
rect -23 258 -19 268
rect -15 258 -11 268
rect -668 172 -663 182
rect -654 172 -649 182
rect -637 172 -632 182
rect -625 172 -621 182
rect -1182 131 -1178 141
rect -1174 131 -1170 141
rect -1149 132 -1145 142
rect -1141 132 -1137 142
rect -1121 133 -1116 143
rect -1107 133 -1102 143
rect -1090 133 -1085 143
rect -1035 133 -1030 143
rect -1021 133 -1016 143
rect -1004 133 -999 143
rect -1065 116 -1061 126
rect -1057 116 -1053 126
rect -979 116 -975 126
rect -971 116 -967 126
rect -949 116 -945 136
rect -930 116 -926 136
rect -911 118 -907 128
rect -903 118 -899 128
rect -604 150 -600 160
rect -596 150 -592 160
rect -296 151 -292 161
rect -288 151 -284 161
rect -263 152 -259 162
rect -255 152 -251 162
rect -235 153 -230 163
rect -221 153 -216 163
rect -204 153 -199 163
rect -149 153 -144 163
rect -135 153 -130 163
rect -118 153 -113 163
rect -179 136 -175 146
rect -171 136 -167 146
rect -93 136 -89 146
rect -85 136 -81 146
rect -63 136 -59 156
rect -44 136 -40 156
rect -25 138 -21 148
rect -17 138 -13 148
rect -989 45 -984 55
rect -975 45 -970 55
rect -958 45 -953 55
rect -667 52 -662 62
rect -653 52 -648 62
rect -636 52 -631 62
rect -933 28 -929 38
rect -925 28 -921 38
rect -611 35 -607 45
rect -603 35 -599 45
rect -574 40 -570 60
rect -555 40 -551 60
rect -536 42 -532 52
rect -528 42 -524 52
rect -296 34 -292 44
rect -288 34 -284 44
rect -263 35 -259 45
rect -255 35 -251 45
rect -235 36 -230 46
rect -221 36 -216 46
rect -204 36 -199 46
rect -149 36 -144 46
rect -135 36 -130 46
rect -118 36 -113 46
rect -179 19 -175 29
rect -171 19 -167 29
rect -93 19 -89 29
rect -85 19 -81 29
rect -63 19 -59 39
rect -44 19 -40 39
rect -25 21 -21 31
rect -17 21 -13 31
<< polysilicon >>
rect -1177 796 -1175 800
rect -1144 797 -1142 801
rect -1113 798 -1110 802
rect -1099 798 -1096 802
rect -1027 798 -1024 802
rect -1013 798 -1010 802
rect -944 791 -942 794
rect -933 791 -931 794
rect -1177 767 -1175 786
rect -1144 768 -1142 787
rect -1113 768 -1110 788
rect -1177 756 -1175 762
rect -1144 757 -1142 763
rect -1113 751 -1110 763
rect -1099 760 -1096 788
rect -1060 781 -1058 785
rect -1099 751 -1096 755
rect -1060 752 -1058 771
rect -1027 768 -1024 788
rect -1027 751 -1024 763
rect -1013 760 -1010 788
rect -974 781 -972 785
rect -906 783 -904 787
rect -1013 751 -1010 755
rect -974 752 -972 771
rect -1060 741 -1058 747
rect -944 747 -942 771
rect -933 747 -931 771
rect -906 754 -904 773
rect -974 741 -972 747
rect -906 743 -904 749
rect -1113 738 -1110 741
rect -1099 738 -1096 741
rect -1027 738 -1024 741
rect -1013 738 -1010 741
rect -944 739 -942 742
rect -933 739 -931 742
rect -981 710 -978 714
rect -967 710 -964 714
rect -981 680 -978 700
rect -981 663 -978 675
rect -967 672 -964 700
rect -928 693 -926 697
rect -967 663 -964 667
rect -928 664 -926 683
rect -928 653 -926 659
rect -981 650 -978 653
rect -967 650 -964 653
rect -638 640 -635 644
rect -624 640 -621 644
rect -638 610 -635 630
rect -638 593 -635 605
rect -624 602 -621 630
rect -585 623 -583 627
rect -624 593 -621 597
rect -585 594 -583 613
rect -1179 584 -1177 588
rect -1146 585 -1144 589
rect -1115 586 -1112 590
rect -1101 586 -1098 590
rect -1029 586 -1026 590
rect -1015 586 -1012 590
rect -585 583 -583 589
rect -946 579 -944 582
rect -935 579 -933 582
rect -638 580 -635 583
rect -624 580 -621 583
rect -1179 555 -1177 574
rect -1146 556 -1144 575
rect -1115 556 -1112 576
rect -1179 544 -1177 550
rect -1146 545 -1144 551
rect -1115 539 -1112 551
rect -1101 548 -1098 576
rect -1062 569 -1060 573
rect -1101 539 -1098 543
rect -1062 540 -1060 559
rect -1029 556 -1026 576
rect -1029 539 -1026 551
rect -1015 548 -1012 576
rect -976 569 -974 573
rect -908 571 -906 575
rect -1015 539 -1012 543
rect -976 540 -974 559
rect -1062 529 -1060 535
rect -946 535 -944 559
rect -935 535 -933 559
rect -908 542 -906 561
rect -512 557 -510 560
rect -501 557 -499 560
rect -490 557 -488 560
rect -480 557 -478 560
rect -642 539 -639 543
rect -628 539 -625 543
rect -613 539 -610 543
rect -976 529 -974 535
rect -908 531 -906 537
rect -1115 526 -1112 529
rect -1101 526 -1098 529
rect -1029 526 -1026 529
rect -1015 526 -1012 529
rect -946 527 -944 530
rect -935 527 -933 530
rect -983 498 -980 502
rect -969 498 -966 502
rect -983 468 -980 488
rect -983 451 -980 463
rect -969 460 -966 488
rect -930 481 -928 485
rect -642 484 -639 529
rect -628 484 -625 529
rect -613 484 -610 529
rect -581 517 -579 521
rect -446 537 -444 541
rect -581 488 -579 507
rect -969 451 -966 455
rect -930 452 -928 471
rect -581 477 -579 483
rect -512 482 -510 517
rect -501 482 -499 517
rect -490 482 -488 517
rect -480 482 -478 517
rect -446 508 -444 527
rect -446 497 -444 503
rect -512 474 -510 477
rect -501 474 -499 477
rect -490 474 -488 477
rect -480 474 -478 477
rect -642 465 -639 469
rect -628 465 -625 469
rect -613 465 -610 469
rect -930 441 -928 447
rect -983 438 -980 441
rect -969 438 -966 441
rect -645 417 -642 421
rect -631 417 -628 421
rect -620 417 -617 421
rect -611 417 -608 421
rect -1180 369 -1178 373
rect -1147 370 -1145 374
rect -1116 371 -1113 375
rect -1102 371 -1099 375
rect -1030 371 -1027 375
rect -1016 371 -1013 375
rect -947 364 -945 367
rect -936 364 -934 367
rect -1180 340 -1178 359
rect -1147 341 -1145 360
rect -1116 341 -1113 361
rect -1180 329 -1178 335
rect -1147 330 -1145 336
rect -1116 324 -1113 336
rect -1102 333 -1099 361
rect -1063 354 -1061 358
rect -1102 324 -1099 328
rect -1063 325 -1061 344
rect -1030 341 -1027 361
rect -1030 324 -1027 336
rect -1016 333 -1013 361
rect -977 354 -975 358
rect -645 362 -642 407
rect -631 362 -628 407
rect -620 373 -617 407
rect -619 368 -617 373
rect -611 368 -608 407
rect -584 395 -582 399
rect -289 398 -287 402
rect -256 399 -254 403
rect -225 400 -222 404
rect -211 400 -208 404
rect -139 400 -136 404
rect -125 400 -122 404
rect -56 393 -54 396
rect -45 393 -43 396
rect -620 362 -617 368
rect -584 366 -582 385
rect -289 369 -287 388
rect -256 370 -254 389
rect -225 370 -222 390
rect -611 362 -608 363
rect -909 356 -907 360
rect -1016 324 -1013 328
rect -977 325 -975 344
rect -1063 314 -1061 320
rect -947 320 -945 344
rect -936 320 -934 344
rect -909 327 -907 346
rect -584 355 -582 361
rect -289 358 -287 364
rect -256 359 -254 365
rect -225 353 -222 365
rect -211 362 -208 390
rect -172 383 -170 387
rect -211 353 -208 357
rect -172 354 -170 373
rect -139 370 -136 390
rect -139 353 -136 365
rect -125 362 -122 390
rect -86 383 -84 387
rect -18 385 -16 389
rect -125 353 -122 357
rect -86 354 -84 373
rect -172 343 -170 349
rect -56 349 -54 373
rect -45 349 -43 373
rect -18 356 -16 375
rect -86 343 -84 349
rect -18 345 -16 351
rect -645 339 -642 342
rect -631 339 -628 342
rect -620 339 -617 342
rect -611 339 -608 342
rect -225 340 -222 343
rect -211 340 -208 343
rect -139 340 -136 343
rect -125 340 -122 343
rect -56 341 -54 344
rect -45 341 -43 344
rect -977 314 -975 320
rect -909 316 -907 322
rect -1116 311 -1113 314
rect -1102 311 -1099 314
rect -1030 311 -1027 314
rect -1016 311 -1013 314
rect -947 312 -945 315
rect -936 312 -934 315
rect -984 283 -981 287
rect -970 283 -967 287
rect -656 283 -653 287
rect -642 283 -639 287
rect -289 281 -287 285
rect -256 282 -254 286
rect -225 283 -222 287
rect -211 283 -208 287
rect -139 283 -136 287
rect -125 283 -122 287
rect -984 253 -981 273
rect -984 236 -981 248
rect -970 245 -967 273
rect -931 266 -929 270
rect -970 236 -967 240
rect -931 237 -929 256
rect -656 253 -653 273
rect -656 236 -653 248
rect -642 245 -639 273
rect -56 276 -54 279
rect -45 276 -43 279
rect -603 266 -601 270
rect -642 236 -639 240
rect -603 237 -601 256
rect -551 254 -549 259
rect -540 254 -538 259
rect -527 254 -525 259
rect -931 226 -929 232
rect -603 226 -601 232
rect -984 223 -981 226
rect -970 223 -967 226
rect -656 223 -653 226
rect -642 223 -639 226
rect -289 252 -287 271
rect -256 253 -254 272
rect -225 253 -222 273
rect -485 243 -483 247
rect -289 241 -287 247
rect -256 242 -254 248
rect -225 236 -222 248
rect -211 245 -208 273
rect -172 266 -170 270
rect -211 236 -208 240
rect -172 237 -170 256
rect -139 253 -136 273
rect -551 189 -549 224
rect -540 189 -538 224
rect -527 189 -525 224
rect -485 214 -483 233
rect -139 236 -136 248
rect -125 245 -122 273
rect -86 266 -84 270
rect -18 268 -16 272
rect -125 236 -122 240
rect -86 237 -84 256
rect -172 226 -170 232
rect -56 232 -54 256
rect -45 232 -43 256
rect -18 239 -16 258
rect -86 226 -84 232
rect -18 228 -16 234
rect -225 223 -222 226
rect -211 223 -208 226
rect -139 223 -136 226
rect -125 223 -122 226
rect -56 224 -54 227
rect -45 224 -43 227
rect -485 203 -483 209
rect -660 182 -657 186
rect -646 182 -643 186
rect -631 182 -628 186
rect -551 182 -549 185
rect -540 182 -538 185
rect -527 182 -525 185
rect -1177 141 -1175 145
rect -1144 142 -1142 146
rect -1113 143 -1110 147
rect -1099 143 -1096 147
rect -1027 143 -1024 147
rect -1013 143 -1010 147
rect -944 136 -942 139
rect -933 136 -931 139
rect -1177 112 -1175 131
rect -1144 113 -1142 132
rect -1113 113 -1110 133
rect -1177 101 -1175 107
rect -1144 102 -1142 108
rect -1113 96 -1110 108
rect -1099 105 -1096 133
rect -1060 126 -1058 130
rect -1099 96 -1096 100
rect -1060 97 -1058 116
rect -1027 113 -1024 133
rect -1027 96 -1024 108
rect -1013 105 -1010 133
rect -974 126 -972 130
rect -906 128 -904 132
rect -660 127 -657 172
rect -646 127 -643 172
rect -631 127 -628 172
rect -599 160 -597 164
rect -291 161 -289 165
rect -258 162 -256 166
rect -227 163 -224 167
rect -213 163 -210 167
rect -141 163 -138 167
rect -127 163 -124 167
rect -58 156 -56 159
rect -47 156 -45 159
rect -599 131 -597 150
rect -291 132 -289 151
rect -258 133 -256 152
rect -227 133 -224 153
rect -1013 96 -1010 100
rect -974 97 -972 116
rect -1060 86 -1058 92
rect -944 92 -942 116
rect -933 92 -931 116
rect -906 99 -904 118
rect -599 120 -597 126
rect -291 121 -289 127
rect -258 122 -256 128
rect -227 116 -224 128
rect -213 125 -210 153
rect -174 146 -172 150
rect -213 116 -210 120
rect -174 117 -172 136
rect -141 133 -138 153
rect -660 108 -657 112
rect -646 108 -643 112
rect -631 108 -628 112
rect -141 116 -138 128
rect -127 125 -124 153
rect -88 146 -86 150
rect -20 148 -18 152
rect -127 116 -124 120
rect -88 117 -86 136
rect -174 106 -172 112
rect -58 112 -56 136
rect -47 112 -45 136
rect -20 119 -18 138
rect -88 106 -86 112
rect -20 108 -18 114
rect -227 103 -224 106
rect -213 103 -210 106
rect -141 103 -138 106
rect -127 103 -124 106
rect -58 104 -56 107
rect -47 104 -45 107
rect -974 86 -972 92
rect -906 88 -904 94
rect -1113 83 -1110 86
rect -1099 83 -1096 86
rect -1027 83 -1024 86
rect -1013 83 -1010 86
rect -944 84 -942 87
rect -933 84 -931 87
rect -659 62 -656 66
rect -645 62 -642 66
rect -981 55 -978 59
rect -967 55 -964 59
rect -569 60 -567 63
rect -558 60 -556 63
rect -981 25 -978 45
rect -981 8 -978 20
rect -967 17 -964 45
rect -928 38 -926 42
rect -659 32 -656 52
rect -967 8 -964 12
rect -928 9 -926 28
rect -659 15 -656 27
rect -645 24 -642 52
rect -606 45 -604 49
rect -531 52 -529 56
rect -291 44 -289 48
rect -258 45 -256 49
rect -227 46 -224 50
rect -213 46 -210 50
rect -141 46 -138 50
rect -127 46 -124 50
rect -645 15 -642 19
rect -606 16 -604 35
rect -569 16 -567 40
rect -558 16 -556 40
rect -531 23 -529 42
rect -58 39 -56 42
rect -47 39 -45 42
rect -531 12 -529 18
rect -291 15 -289 34
rect -258 16 -256 35
rect -227 16 -224 36
rect -606 5 -604 11
rect -569 8 -567 11
rect -558 8 -556 11
rect -928 -2 -926 4
rect -659 2 -656 5
rect -645 2 -642 5
rect -291 4 -289 10
rect -258 5 -256 11
rect -227 -1 -224 11
rect -213 8 -210 36
rect -174 29 -172 33
rect -213 -1 -210 3
rect -174 0 -172 19
rect -141 16 -138 36
rect -981 -5 -978 -2
rect -967 -5 -964 -2
rect -141 -1 -138 11
rect -127 8 -124 36
rect -88 29 -86 33
rect -20 31 -18 35
rect -127 -1 -124 3
rect -88 0 -86 19
rect -174 -11 -172 -5
rect -58 -5 -56 19
rect -47 -5 -45 19
rect -20 2 -18 21
rect -88 -11 -86 -5
rect -20 -9 -18 -3
rect -227 -14 -224 -11
rect -213 -14 -210 -11
rect -141 -14 -138 -11
rect -127 -14 -124 -11
rect -58 -13 -56 -10
rect -47 -13 -45 -10
<< polycontact >>
rect -1181 770 -1177 774
rect -1148 771 -1144 775
rect -1115 763 -1110 768
rect -1101 755 -1096 760
rect -1064 755 -1060 759
rect -1029 763 -1024 768
rect -1015 755 -1010 760
rect -978 755 -974 759
rect -948 758 -944 762
rect -937 758 -933 762
rect -910 757 -906 761
rect -983 675 -978 680
rect -969 667 -964 672
rect -932 667 -928 671
rect -640 605 -635 610
rect -626 597 -621 602
rect -589 597 -585 601
rect -1183 558 -1179 562
rect -1150 559 -1146 563
rect -1117 551 -1112 556
rect -1103 543 -1098 548
rect -1066 543 -1062 547
rect -1031 551 -1026 556
rect -1017 543 -1012 548
rect -980 543 -976 547
rect -950 546 -946 550
rect -939 546 -935 550
rect -912 545 -908 549
rect -647 504 -642 509
rect -985 463 -980 468
rect -633 496 -628 501
rect -618 487 -613 492
rect -585 491 -581 495
rect -516 505 -512 509
rect -971 455 -966 460
rect -934 455 -930 459
rect -505 498 -501 502
rect -494 491 -490 495
rect -484 492 -480 496
rect -450 511 -446 515
rect -650 382 -645 387
rect -1184 343 -1180 347
rect -1151 344 -1147 348
rect -1118 336 -1113 341
rect -1104 328 -1099 333
rect -1067 328 -1063 332
rect -1032 336 -1027 341
rect -636 374 -631 379
rect -624 368 -619 373
rect -588 369 -584 373
rect -613 363 -608 368
rect -293 372 -289 376
rect -260 373 -256 377
rect -1018 328 -1013 333
rect -981 328 -977 332
rect -951 331 -947 335
rect -940 331 -936 335
rect -913 330 -909 334
rect -227 365 -222 370
rect -213 357 -208 362
rect -176 357 -172 361
rect -141 365 -136 370
rect -127 357 -122 362
rect -90 357 -86 361
rect -60 360 -56 364
rect -49 360 -45 364
rect -22 359 -18 363
rect -986 248 -981 253
rect -972 240 -967 245
rect -935 240 -931 244
rect -658 248 -653 253
rect -644 240 -639 245
rect -607 240 -603 244
rect -293 255 -289 259
rect -260 256 -256 260
rect -227 248 -222 253
rect -213 240 -208 245
rect -176 240 -172 244
rect -141 248 -136 253
rect -555 211 -551 215
rect -544 205 -540 209
rect -531 198 -527 202
rect -489 217 -485 221
rect -127 240 -122 245
rect -90 240 -86 244
rect -60 243 -56 247
rect -49 243 -45 247
rect -22 242 -18 246
rect -665 147 -660 152
rect -1181 115 -1177 119
rect -1148 116 -1144 120
rect -1115 108 -1110 113
rect -1101 100 -1096 105
rect -1064 100 -1060 104
rect -1029 108 -1024 113
rect -651 139 -646 144
rect -636 130 -631 135
rect -603 134 -599 138
rect -295 135 -291 139
rect -262 136 -258 140
rect -1015 100 -1010 105
rect -978 100 -974 104
rect -948 103 -944 107
rect -937 103 -933 107
rect -910 102 -906 106
rect -229 128 -224 133
rect -215 120 -210 125
rect -178 120 -174 124
rect -143 128 -138 133
rect -129 120 -124 125
rect -92 120 -88 124
rect -62 123 -58 127
rect -51 123 -47 127
rect -24 122 -20 126
rect -983 20 -978 25
rect -969 12 -964 17
rect -932 12 -928 16
rect -661 27 -656 32
rect -647 19 -642 24
rect -610 19 -606 23
rect -573 27 -569 31
rect -562 27 -558 31
rect -535 26 -531 30
rect -295 18 -291 22
rect -262 19 -258 23
rect -229 11 -224 16
rect -215 3 -210 8
rect -178 3 -174 7
rect -143 11 -138 16
rect -129 3 -124 8
rect -92 3 -88 7
rect -62 6 -58 10
rect -51 6 -47 10
rect -24 5 -20 9
<< metal1 >>
rect -1189 802 -1164 806
rect -1156 803 -1131 807
rect -1121 806 -1052 810
rect -1035 806 -966 810
rect -1182 796 -1178 802
rect -1149 797 -1145 803
rect -1121 798 -1116 806
rect -1090 798 -1085 806
rect -1058 791 -1053 806
rect -1035 798 -1030 806
rect -1004 798 -999 806
rect -1174 774 -1170 786
rect -1141 775 -1137 787
rect -1189 770 -1181 774
rect -1174 770 -1162 774
rect -1156 771 -1148 775
rect -1141 771 -1129 775
rect -1174 767 -1170 770
rect -1141 768 -1137 771
rect -1107 768 -1102 788
rect -1072 787 -1047 791
rect -972 791 -967 806
rect -955 797 -906 801
rect -949 791 -945 797
rect -912 793 -906 797
rect -1065 781 -1061 787
rect -1118 763 -1115 768
rect -1107 764 -1085 768
rect -1182 753 -1178 762
rect -1149 754 -1145 763
rect -1118 755 -1101 760
rect -1090 759 -1085 764
rect -1057 759 -1053 771
rect -1021 768 -1016 788
rect -986 787 -961 791
rect -979 781 -975 787
rect -915 789 -893 793
rect -911 783 -907 789
rect -1032 763 -1029 768
rect -1021 764 -999 768
rect -1090 755 -1064 759
rect -1057 755 -1045 759
rect -1032 755 -1015 760
rect -1004 759 -999 764
rect -971 759 -967 771
rect -1004 755 -978 759
rect -971 755 -959 759
rect -930 761 -926 771
rect -903 761 -899 773
rect -930 757 -910 761
rect -903 757 -891 761
rect -1186 749 -1166 753
rect -1153 750 -1133 754
rect -1090 751 -1085 755
rect -1057 752 -1053 755
rect -1004 751 -999 755
rect -971 752 -967 755
rect -930 754 -926 757
rect -903 754 -899 757
rect -1121 737 -1116 741
rect -1065 738 -1061 747
rect -940 751 -926 754
rect -940 747 -936 751
rect -1069 737 -1049 738
rect -1121 734 -1049 737
rect -1035 737 -1030 741
rect -979 738 -975 747
rect -983 737 -963 738
rect -1035 734 -963 737
rect -949 736 -945 742
rect -930 740 -926 742
rect -911 740 -907 749
rect -930 736 -895 740
rect -1121 733 -1085 734
rect -1035 733 -999 734
rect -949 733 -926 736
rect -989 718 -920 722
rect -989 710 -984 718
rect -958 710 -953 718
rect -926 703 -921 718
rect -975 680 -970 700
rect -940 699 -915 703
rect -933 693 -929 699
rect -986 675 -983 680
rect -975 676 -953 680
rect -986 667 -969 672
rect -958 671 -953 676
rect -925 671 -921 683
rect -958 667 -932 671
rect -925 667 -913 671
rect -958 663 -953 667
rect -925 664 -921 667
rect -989 649 -984 653
rect -933 650 -929 659
rect -937 649 -917 650
rect -989 646 -917 649
rect -646 648 -577 652
rect -989 645 -953 646
rect -646 640 -641 648
rect -615 640 -610 648
rect -583 633 -578 648
rect -632 610 -627 630
rect -597 629 -572 633
rect -590 623 -586 629
rect -643 605 -640 610
rect -632 606 -610 610
rect -1191 590 -1166 594
rect -1158 591 -1133 595
rect -1123 594 -1054 598
rect -1037 594 -968 598
rect -643 597 -626 602
rect -615 601 -610 606
rect -582 601 -578 613
rect -615 597 -589 601
rect -582 597 -549 601
rect -1184 584 -1180 590
rect -1151 585 -1147 591
rect -1123 586 -1118 594
rect -1092 586 -1087 594
rect -1060 579 -1055 594
rect -1037 586 -1032 594
rect -1006 586 -1001 594
rect -1176 562 -1172 574
rect -1143 563 -1139 575
rect -1191 558 -1183 562
rect -1176 558 -1164 562
rect -1158 559 -1150 563
rect -1143 559 -1131 563
rect -1176 555 -1172 558
rect -1143 556 -1139 559
rect -1109 556 -1104 576
rect -1074 575 -1049 579
rect -974 579 -969 594
rect -615 593 -610 597
rect -582 594 -578 597
rect -957 585 -908 589
rect -951 579 -947 585
rect -914 581 -908 585
rect -1067 569 -1063 575
rect -1120 551 -1117 556
rect -1109 552 -1087 556
rect -1184 541 -1180 550
rect -1151 542 -1147 551
rect -1120 543 -1103 548
rect -1092 547 -1087 552
rect -1059 547 -1055 559
rect -1023 556 -1018 576
rect -988 575 -963 579
rect -981 569 -977 575
rect -917 577 -895 581
rect -646 579 -641 583
rect -590 580 -586 589
rect -594 579 -574 580
rect -913 571 -909 577
rect -646 576 -574 579
rect -646 575 -610 576
rect -1034 551 -1031 556
rect -1023 552 -1001 556
rect -1092 543 -1066 547
rect -1059 543 -1047 547
rect -1034 543 -1017 548
rect -1006 547 -1001 552
rect -973 547 -969 559
rect -1006 543 -980 547
rect -973 543 -961 547
rect -932 549 -928 559
rect -905 549 -901 561
rect -932 545 -912 549
rect -905 545 -893 549
rect -650 547 -578 551
rect -1188 537 -1168 541
rect -1155 538 -1135 542
rect -1092 539 -1087 543
rect -1059 540 -1055 543
rect -1006 539 -1001 543
rect -973 540 -969 543
rect -932 542 -928 545
rect -905 542 -901 545
rect -1123 525 -1118 529
rect -1067 526 -1063 535
rect -942 539 -928 542
rect -942 535 -938 539
rect -650 539 -645 547
rect -619 539 -614 547
rect -1071 525 -1051 526
rect -1123 522 -1051 525
rect -1037 525 -1032 529
rect -981 526 -977 535
rect -985 525 -965 526
rect -1037 522 -965 525
rect -951 524 -947 530
rect -932 528 -928 530
rect -913 528 -909 537
rect -584 531 -579 547
rect -932 524 -897 528
rect -1123 521 -1087 522
rect -1037 521 -1001 522
rect -951 521 -928 524
rect -991 506 -922 510
rect -636 509 -631 529
rect -607 509 -603 529
rect -593 527 -568 531
rect -991 498 -986 506
rect -960 498 -955 506
rect -928 491 -923 506
rect -636 505 -603 509
rect -586 517 -582 527
rect -607 495 -603 505
rect -578 495 -574 507
rect -552 509 -549 597
rect -517 563 -448 567
rect -517 557 -513 563
rect -455 547 -448 563
rect -455 543 -433 547
rect -451 537 -447 543
rect -552 505 -516 509
rect -477 508 -471 517
rect -443 515 -439 527
rect -458 511 -450 515
rect -443 511 -431 515
rect -458 508 -454 511
rect -443 508 -439 511
rect -477 504 -454 508
rect -548 498 -505 502
rect -548 495 -545 498
rect -977 468 -972 488
rect -942 487 -917 491
rect -607 491 -585 495
rect -578 491 -545 495
rect -538 491 -494 495
rect -935 481 -931 487
rect -607 484 -603 491
rect -578 488 -574 491
rect -988 463 -985 468
rect -977 464 -955 468
rect -988 455 -971 460
rect -960 459 -955 464
rect -927 459 -923 471
rect -586 474 -582 483
rect -590 470 -570 474
rect -650 461 -646 469
rect -590 461 -585 470
rect -960 455 -934 459
rect -927 455 -915 459
rect -650 456 -585 461
rect -960 451 -955 455
rect -927 452 -923 455
rect -991 437 -986 441
rect -935 438 -931 447
rect -939 437 -919 438
rect -991 434 -919 437
rect -991 433 -955 434
rect -653 425 -581 429
rect -653 417 -648 425
rect -626 417 -622 425
rect -606 417 -602 425
rect -587 409 -582 425
rect -639 387 -634 407
rect -616 387 -612 407
rect -596 405 -571 409
rect -589 395 -585 405
rect -1192 375 -1167 379
rect -1159 376 -1134 380
rect -1124 379 -1055 383
rect -1038 379 -969 383
rect -639 383 -601 387
rect -1185 369 -1181 375
rect -1152 370 -1148 376
rect -1124 371 -1119 379
rect -1093 371 -1088 379
rect -1061 364 -1056 379
rect -1038 371 -1033 379
rect -1007 371 -1002 379
rect -1177 347 -1173 359
rect -1144 348 -1140 360
rect -1192 343 -1184 347
rect -1177 343 -1165 347
rect -1159 344 -1151 348
rect -1144 344 -1132 348
rect -1177 340 -1173 343
rect -1144 341 -1140 344
rect -1110 341 -1105 361
rect -1075 360 -1050 364
rect -975 364 -970 379
rect -958 370 -909 374
rect -605 373 -601 383
rect -581 373 -577 385
rect -538 373 -533 491
rect -477 488 -471 504
rect -507 485 -471 488
rect -507 482 -503 485
rect -486 482 -482 485
rect -517 473 -513 477
rect -495 473 -491 477
rect -477 473 -471 477
rect -451 473 -447 503
rect -517 470 -447 473
rect -301 404 -276 408
rect -268 405 -243 409
rect -233 408 -164 412
rect -147 408 -78 412
rect -294 398 -290 404
rect -261 399 -257 405
rect -233 400 -228 408
rect -202 400 -197 408
rect -170 393 -165 408
rect -147 400 -142 408
rect -116 400 -111 408
rect -286 376 -282 388
rect -253 377 -249 389
rect -952 364 -948 370
rect -915 366 -909 370
rect -605 369 -588 373
rect -581 369 -533 373
rect -301 372 -293 376
rect -286 372 -274 376
rect -268 373 -260 377
rect -253 373 -241 377
rect -286 369 -282 372
rect -253 370 -249 373
rect -219 370 -214 390
rect -184 389 -159 393
rect -84 393 -79 408
rect -67 399 -18 403
rect -61 393 -57 399
rect -24 395 -18 399
rect -177 383 -173 389
rect -1068 354 -1064 360
rect -1121 336 -1118 341
rect -1110 337 -1088 341
rect -1185 326 -1181 335
rect -1152 327 -1148 336
rect -1121 328 -1104 333
rect -1093 332 -1088 337
rect -1060 332 -1056 344
rect -1024 341 -1019 361
rect -989 360 -964 364
rect -982 354 -978 360
rect -918 362 -896 366
rect -605 362 -601 369
rect -581 366 -577 369
rect -914 356 -910 362
rect -1035 336 -1032 341
rect -1024 337 -1002 341
rect -1093 328 -1067 332
rect -1060 328 -1048 332
rect -1035 328 -1018 333
rect -1007 332 -1002 337
rect -974 332 -970 344
rect -1007 328 -981 332
rect -974 328 -962 332
rect -933 334 -929 344
rect -906 334 -902 346
rect -230 365 -227 370
rect -219 366 -197 370
rect -589 352 -585 361
rect -294 355 -290 364
rect -261 356 -257 365
rect -230 357 -213 362
rect -202 361 -197 366
rect -169 361 -165 373
rect -133 370 -128 390
rect -98 389 -73 393
rect -91 383 -87 389
rect -27 391 -5 395
rect -23 385 -19 391
rect -144 365 -141 370
rect -133 366 -111 370
rect -202 357 -176 361
rect -169 357 -157 361
rect -144 357 -127 362
rect -116 361 -111 366
rect -83 361 -79 373
rect -116 357 -90 361
rect -83 357 -71 361
rect -42 363 -38 373
rect -15 363 -11 375
rect -42 359 -22 363
rect -15 359 -3 363
rect -593 348 -573 352
rect -298 351 -278 355
rect -265 352 -245 356
rect -202 353 -197 357
rect -169 354 -165 357
rect -653 338 -649 342
rect -593 338 -588 348
rect -653 334 -588 338
rect -116 353 -111 357
rect -83 354 -79 357
rect -42 356 -38 359
rect -15 356 -11 359
rect -233 339 -228 343
rect -177 340 -173 349
rect -52 353 -38 356
rect -52 349 -48 353
rect -181 339 -161 340
rect -233 336 -161 339
rect -147 339 -142 343
rect -91 340 -87 349
rect -95 339 -75 340
rect -147 336 -75 339
rect -61 338 -57 344
rect -42 342 -38 344
rect -23 342 -19 351
rect -42 338 -7 342
rect -233 335 -197 336
rect -147 335 -111 336
rect -61 335 -38 338
rect -933 330 -913 334
rect -906 330 -894 334
rect -1189 322 -1169 326
rect -1156 323 -1136 327
rect -1093 324 -1088 328
rect -1060 325 -1056 328
rect -1007 324 -1002 328
rect -974 325 -970 328
rect -933 327 -929 330
rect -906 327 -902 330
rect -1124 310 -1119 314
rect -1068 311 -1064 320
rect -943 324 -929 327
rect -943 320 -939 324
rect -1072 310 -1052 311
rect -1124 307 -1052 310
rect -1038 310 -1033 314
rect -982 311 -978 320
rect -986 310 -966 311
rect -1038 307 -966 310
rect -952 309 -948 315
rect -933 313 -929 315
rect -914 313 -910 322
rect -933 309 -898 313
rect -1124 306 -1088 307
rect -1038 306 -1002 307
rect -952 306 -929 309
rect -992 291 -923 295
rect -664 291 -595 295
rect -992 283 -987 291
rect -961 283 -956 291
rect -929 276 -924 291
rect -664 283 -659 291
rect -633 283 -628 291
rect -978 253 -973 273
rect -943 272 -918 276
rect -601 276 -596 291
rect -301 287 -276 291
rect -268 288 -243 292
rect -233 291 -164 295
rect -147 291 -78 295
rect -294 281 -290 287
rect -261 282 -257 288
rect -233 283 -228 291
rect -202 283 -197 291
rect -936 266 -932 272
rect -989 248 -986 253
rect -978 249 -956 253
rect -989 240 -972 245
rect -961 244 -956 249
rect -928 244 -924 256
rect -650 253 -645 273
rect -615 272 -590 276
rect -608 266 -604 272
rect -170 276 -165 291
rect -147 283 -142 291
rect -116 283 -111 291
rect -562 262 -486 266
rect -661 248 -658 253
rect -650 249 -628 253
rect -961 240 -935 244
rect -928 240 -916 244
rect -661 240 -644 245
rect -633 244 -628 249
rect -600 244 -596 256
rect -556 254 -552 262
rect -633 240 -607 244
rect -600 240 -581 244
rect -961 236 -956 240
rect -928 237 -924 240
rect -633 236 -628 240
rect -600 237 -596 240
rect -992 222 -987 226
rect -936 223 -932 232
rect -940 222 -920 223
rect -992 219 -920 222
rect -664 222 -659 226
rect -608 223 -604 232
rect -612 222 -592 223
rect -664 219 -592 222
rect -992 218 -956 219
rect -664 218 -628 219
rect -585 215 -581 240
rect -494 253 -487 262
rect -286 259 -282 271
rect -253 260 -249 272
rect -301 255 -293 259
rect -286 255 -274 259
rect -268 256 -260 260
rect -253 256 -241 260
rect -494 249 -472 253
rect -286 252 -282 255
rect -253 253 -249 256
rect -219 253 -214 273
rect -184 272 -159 276
rect -84 276 -79 291
rect -67 282 -18 286
rect -61 276 -57 282
rect -24 278 -18 282
rect -177 266 -173 272
rect -490 243 -486 249
rect -230 248 -227 253
rect -219 249 -197 253
rect -294 238 -290 247
rect -261 239 -257 248
rect -230 240 -213 245
rect -202 244 -197 249
rect -169 244 -165 256
rect -133 253 -128 273
rect -98 272 -73 276
rect -91 266 -87 272
rect -27 274 -5 278
rect -23 268 -19 274
rect -144 248 -141 253
rect -133 249 -111 253
rect -202 240 -176 244
rect -169 240 -157 244
rect -144 240 -127 245
rect -116 244 -111 249
rect -83 244 -79 256
rect -116 240 -90 244
rect -83 240 -71 244
rect -42 246 -38 256
rect -15 246 -11 258
rect -42 242 -22 246
rect -15 242 -3 246
rect -298 234 -278 238
rect -265 235 -245 239
rect -202 236 -197 240
rect -169 237 -165 240
rect -585 211 -555 215
rect -516 214 -510 224
rect -482 221 -478 233
rect -116 236 -111 240
rect -83 237 -79 240
rect -42 239 -38 242
rect -15 239 -11 242
rect -233 222 -228 226
rect -177 223 -173 232
rect -52 236 -38 239
rect -52 232 -48 236
rect -181 222 -161 223
rect -497 217 -489 221
rect -482 217 -470 221
rect -233 219 -161 222
rect -147 222 -142 226
rect -91 223 -87 232
rect -95 222 -75 223
rect -147 219 -75 222
rect -61 221 -57 227
rect -42 225 -38 227
rect -23 225 -19 234
rect -42 221 -7 225
rect -233 218 -197 219
rect -147 218 -111 219
rect -61 218 -38 221
rect -497 214 -493 217
rect -482 214 -478 217
rect -516 210 -493 214
rect -568 198 -531 202
rect -668 190 -596 194
rect -668 182 -663 190
rect -637 182 -632 190
rect -602 174 -597 190
rect -1189 147 -1164 151
rect -1156 148 -1131 152
rect -1121 151 -1052 155
rect -1035 151 -966 155
rect -654 152 -649 172
rect -625 152 -621 172
rect -611 170 -586 174
rect -1182 141 -1178 147
rect -1149 142 -1145 148
rect -1121 143 -1116 151
rect -1090 143 -1085 151
rect -1058 136 -1053 151
rect -1035 143 -1030 151
rect -1004 143 -999 151
rect -1174 119 -1170 131
rect -1141 120 -1137 132
rect -1189 115 -1181 119
rect -1174 115 -1162 119
rect -1156 116 -1148 120
rect -1141 116 -1129 120
rect -1174 112 -1170 115
rect -1141 113 -1137 116
rect -1107 113 -1102 133
rect -1072 132 -1047 136
rect -972 136 -967 151
rect -654 148 -621 152
rect -604 160 -600 170
rect -955 142 -906 146
rect -949 136 -945 142
rect -912 138 -906 142
rect -625 138 -621 148
rect -596 138 -592 150
rect -568 138 -565 198
rect -516 195 -510 210
rect -546 192 -510 195
rect -546 189 -542 192
rect -516 189 -510 192
rect -556 179 -552 185
rect -534 179 -530 185
rect -490 179 -486 209
rect -556 176 -486 179
rect -303 167 -278 171
rect -270 168 -245 172
rect -235 171 -166 175
rect -149 171 -80 175
rect -296 161 -292 167
rect -263 162 -259 168
rect -235 163 -230 171
rect -204 163 -199 171
rect -172 156 -167 171
rect -149 163 -144 171
rect -118 163 -113 171
rect -288 139 -284 151
rect -255 140 -251 152
rect -1065 126 -1061 132
rect -1118 108 -1115 113
rect -1107 109 -1085 113
rect -1182 98 -1178 107
rect -1149 99 -1145 108
rect -1118 100 -1101 105
rect -1090 104 -1085 109
rect -1057 104 -1053 116
rect -1021 113 -1016 133
rect -986 132 -961 136
rect -979 126 -975 132
rect -915 134 -893 138
rect -911 128 -907 134
rect -708 130 -636 135
rect -625 134 -603 138
rect -596 134 -565 138
rect -303 135 -295 139
rect -288 135 -276 139
rect -270 136 -262 140
rect -255 136 -243 140
rect -1032 108 -1029 113
rect -1021 109 -999 113
rect -1090 100 -1064 104
rect -1057 100 -1045 104
rect -1032 100 -1015 105
rect -1004 104 -999 109
rect -971 104 -967 116
rect -1004 100 -978 104
rect -971 100 -959 104
rect -930 106 -926 116
rect -903 106 -899 118
rect -930 102 -910 106
rect -903 102 -891 106
rect -1186 94 -1166 98
rect -1153 95 -1133 99
rect -1090 96 -1085 100
rect -1057 97 -1053 100
rect -1004 96 -999 100
rect -971 97 -967 100
rect -930 99 -926 102
rect -903 99 -899 102
rect -1121 82 -1116 86
rect -1065 83 -1061 92
rect -940 96 -926 99
rect -940 92 -936 96
rect -1069 82 -1049 83
rect -1121 79 -1049 82
rect -1035 82 -1030 86
rect -979 83 -975 92
rect -983 82 -963 83
rect -1035 79 -963 82
rect -949 81 -945 87
rect -930 85 -926 87
rect -911 85 -907 94
rect -930 81 -895 85
rect -1121 78 -1085 79
rect -1035 78 -999 79
rect -949 78 -926 81
rect -989 63 -920 67
rect -989 55 -984 63
rect -958 55 -953 63
rect -926 48 -921 63
rect -975 25 -970 45
rect -940 44 -915 48
rect -933 38 -929 44
rect -986 20 -983 25
rect -975 21 -953 25
rect -986 12 -969 17
rect -958 16 -953 21
rect -925 16 -921 28
rect -708 16 -702 130
rect -625 127 -621 134
rect -596 131 -592 134
rect -288 132 -284 135
rect -255 133 -251 136
rect -221 133 -216 153
rect -186 152 -161 156
rect -86 156 -81 171
rect -69 162 -20 166
rect -63 156 -59 162
rect -26 158 -20 162
rect -179 146 -175 152
rect -232 128 -229 133
rect -221 129 -199 133
rect -604 117 -600 126
rect -296 118 -292 127
rect -263 119 -259 128
rect -232 120 -215 125
rect -204 124 -199 129
rect -171 124 -167 136
rect -135 133 -130 153
rect -100 152 -75 156
rect -93 146 -89 152
rect -29 154 -7 158
rect -25 148 -21 154
rect -146 128 -143 133
rect -135 129 -113 133
rect -204 120 -178 124
rect -171 120 -159 124
rect -146 120 -129 125
rect -118 124 -113 129
rect -85 124 -81 136
rect -118 120 -92 124
rect -85 120 -73 124
rect -44 126 -40 136
rect -17 126 -13 138
rect -44 122 -24 126
rect -17 122 -5 126
rect -608 113 -588 117
rect -300 114 -280 118
rect -267 115 -247 119
rect -204 116 -199 120
rect -171 117 -167 120
rect -668 104 -664 112
rect -608 104 -603 113
rect -668 99 -603 104
rect -118 116 -113 120
rect -85 117 -81 120
rect -44 119 -40 122
rect -17 119 -13 122
rect -235 102 -230 106
rect -179 103 -175 112
rect -54 116 -40 119
rect -54 112 -50 116
rect -183 102 -163 103
rect -235 99 -163 102
rect -149 102 -144 106
rect -93 103 -89 112
rect -97 102 -77 103
rect -149 99 -77 102
rect -63 101 -59 107
rect -44 105 -40 107
rect -25 105 -21 114
rect -44 101 -9 105
rect -235 98 -199 99
rect -149 98 -113 99
rect -63 98 -40 101
rect -667 70 -598 74
rect -667 62 -662 70
rect -636 62 -631 70
rect -604 55 -599 70
rect -580 66 -531 70
rect -574 60 -570 66
rect -537 62 -531 66
rect -653 32 -648 52
rect -618 51 -593 55
rect -611 45 -607 51
rect -540 58 -518 62
rect -536 52 -532 58
rect -303 50 -278 54
rect -270 51 -245 55
rect -235 54 -166 58
rect -149 54 -80 58
rect -664 27 -661 32
rect -653 28 -631 32
rect -664 22 -647 24
rect -689 19 -647 22
rect -636 23 -631 28
rect -603 23 -599 35
rect -585 27 -573 31
rect -555 30 -551 40
rect -528 30 -524 42
rect -296 44 -292 50
rect -263 45 -259 51
rect -235 46 -230 54
rect -204 46 -199 54
rect -172 39 -167 54
rect -149 46 -144 54
rect -118 46 -113 54
rect -585 23 -582 27
rect -555 26 -535 30
rect -528 26 -516 30
rect -555 23 -551 26
rect -528 23 -524 26
rect -636 19 -610 23
rect -603 19 -582 23
rect -565 20 -551 23
rect -689 16 -686 19
rect -958 12 -932 16
rect -925 12 -686 16
rect -636 15 -631 19
rect -603 16 -599 19
rect -565 16 -561 20
rect -288 22 -284 34
rect -255 23 -251 35
rect -303 18 -295 22
rect -288 18 -276 22
rect -270 19 -262 23
rect -255 19 -243 23
rect -958 8 -953 12
rect -925 9 -921 12
rect -989 -6 -984 -2
rect -933 -5 -929 4
rect -667 1 -662 5
rect -611 2 -607 11
rect -574 5 -570 11
rect -555 9 -551 11
rect -536 9 -532 18
rect -288 15 -284 18
rect -255 16 -251 19
rect -221 16 -216 36
rect -186 35 -161 39
rect -86 39 -81 54
rect -69 45 -20 49
rect -63 39 -59 45
rect -26 41 -20 45
rect -179 29 -175 35
rect -232 11 -229 16
rect -221 12 -199 16
rect -555 5 -520 9
rect -574 2 -551 5
rect -615 1 -595 2
rect -296 1 -292 10
rect -263 2 -259 11
rect -232 3 -215 8
rect -204 7 -199 12
rect -171 7 -167 19
rect -135 16 -130 36
rect -100 35 -75 39
rect -93 29 -89 35
rect -29 37 -7 41
rect -25 31 -21 37
rect -146 11 -143 16
rect -135 12 -113 16
rect -204 3 -178 7
rect -171 3 -159 7
rect -146 3 -129 8
rect -118 7 -113 12
rect -85 7 -81 19
rect -118 3 -92 7
rect -85 3 -73 7
rect -44 9 -40 19
rect -17 9 -13 21
rect -44 5 -24 9
rect -17 5 -5 9
rect -667 -2 -595 1
rect -667 -3 -631 -2
rect -300 -3 -280 1
rect -267 -2 -247 2
rect -204 -1 -199 3
rect -171 0 -167 3
rect -937 -6 -917 -5
rect -989 -9 -917 -6
rect -989 -10 -953 -9
rect -118 -1 -113 3
rect -85 0 -81 3
rect -44 2 -40 5
rect -17 2 -13 5
rect -235 -15 -230 -11
rect -179 -14 -175 -5
rect -54 -1 -40 2
rect -54 -5 -50 -1
rect -183 -15 -163 -14
rect -235 -18 -163 -15
rect -149 -15 -144 -11
rect -93 -14 -89 -5
rect -97 -15 -77 -14
rect -149 -18 -77 -15
rect -63 -16 -59 -10
rect -44 -12 -40 -10
rect -25 -12 -21 -3
rect -44 -16 -9 -12
rect -235 -19 -199 -18
rect -149 -19 -113 -18
rect -63 -19 -40 -16
<< labels >>
rlabel pdcontact -609 40 -609 40 1 vdd
rlabel ndcontact -609 13 -609 13 1 gnd
rlabel metal1 -607 0 -607 0 1 gnd
rlabel metal1 -651 72 -651 72 5 vdd
rlabel ndcontact -665 13 -665 13 1 gnd
rlabel pdcontact -665 57 -665 57 1 vdd
rlabel pdcontact -634 56 -634 56 1 vdd
rlabel polycontact -658 29 -658 29 1 p1
rlabel polycontact -644 21 -644 21 1 g0
rlabel ndiffusion -651 10 -651 10 1 n29
rlabel metal1 -594 21 -594 21 7 p1g0
rlabel ndcontact -601 13 -601 13 1 p1g0
rlabel pdcontact -601 40 -601 40 1 p1g0
rlabel polycontact -608 21 -608 21 1 nand17
rlabel ndcontact -634 10 -634 10 1 nand17
rlabel pdcontact -651 57 -651 57 1 nand17
rlabel pdcontact -534 47 -534 47 1 vdd
rlabel ndcontact -534 20 -534 20 1 gnd
rlabel metal1 -563 3 -563 3 1 gnd
rlabel metal1 -563 68 -563 68 5 vdd
rlabel pdcontact -572 50 -572 50 1 vdd
rlabel ndcontact -554 13 -554 13 1 gnd
rlabel ndcontact -572 14 -572 14 1 gnd
rlabel polycontact -533 28 -533 28 1 nor9
rlabel pdcontact -553 50 -553 50 1 nor9
rlabel ndcontact -563 13 -563 13 1 nor9
rlabel pdiffusion -563 51 -563 51 1 n30
rlabel polycontact -571 29 -571 29 1 p1g0
rlabel polycontact -560 29 -560 29 1 g1
rlabel metal1 -519 28 -519 28 7 c2
rlabel ndcontact -526 20 -526 20 1 c2
rlabel pdcontact -526 47 -526 47 1 c2
rlabel metal1 -652 192 -652 192 5 vdd
rlabel pdcontact -666 177 -666 177 1 vdd
rlabel pdcontact -635 177 -635 177 1 vdd
rlabel ndcontact -666 119 -666 119 1 gnd
rlabel pdcontact -602 155 -602 155 1 vdd
rlabel ndcontact -602 128 -602 128 1 gnd
rlabel metal1 -600 115 -600 115 1 gnd
rlabel pdcontact -606 261 -606 261 1 vdd
rlabel ndcontact -606 234 -606 234 1 gnd
rlabel metal1 -604 221 -604 221 1 gnd
rlabel metal1 -648 293 -648 293 5 vdd
rlabel ndcontact -662 234 -662 234 1 gnd
rlabel pdcontact -662 278 -662 278 1 vdd
rlabel pdcontact -631 277 -631 277 1 vdd
rlabel metal1 -540 264 -540 264 5 vdd
rlabel pdcontact -554 239 -554 239 1 vdd
rlabel pdcontact -488 238 -488 238 1 vdd
rlabel ndcontact -488 211 -488 211 1 gnd
rlabel ndcontact -554 187 -554 187 1 gnd
rlabel ndcontact -532 187 -532 187 1 gnd
rlabel metal1 -519 177 -519 177 1 gnd
rlabel metal1 -637 427 -637 427 5 vdd
rlabel pdcontact -651 412 -651 412 1 vdd
rlabel ndcontact -651 354 -651 354 1 gnd
rlabel pdcontact -587 390 -587 390 1 vdd
rlabel ndcontact -587 363 -587 363 1 gnd
rlabel metal1 -585 350 -585 350 1 gnd
rlabel pdcontact -624 411 -624 411 1 vdd
rlabel pdcontact -604 412 -604 412 1 vdd
rlabel metal1 -634 549 -634 549 5 vdd
rlabel pdcontact -648 534 -648 534 1 vdd
rlabel pdcontact -617 534 -617 534 1 vdd
rlabel ndcontact -648 476 -648 476 1 gnd
rlabel pdcontact -584 512 -584 512 1 vdd
rlabel ndcontact -584 485 -584 485 1 gnd
rlabel metal1 -582 472 -582 472 1 gnd
rlabel pdcontact -588 618 -588 618 1 vdd
rlabel ndcontact -588 591 -588 591 1 gnd
rlabel metal1 -586 578 -586 578 1 gnd
rlabel metal1 -630 650 -630 650 5 vdd
rlabel ndcontact -644 591 -644 591 1 gnd
rlabel pdcontact -644 635 -644 635 1 vdd
rlabel pdcontact -613 634 -613 634 1 vdd
rlabel pdcontact -515 533 -515 533 1 vdd
rlabel pdcontact -449 532 -449 532 1 vdd
rlabel ndcontact -449 505 -449 505 1 gnd
rlabel ndcontact -515 481 -515 481 1 gnd
rlabel ndcontact -493 481 -493 481 1 gnd
rlabel metal1 -480 471 -480 471 1 gnd
rlabel ndcontact -474 481 -474 481 1 gnd
rlabel metal1 -473 565 -473 565 5 vdd
rlabel polycontact -662 149 -662 149 1 p2
rlabel polycontact -649 141 -649 141 1 p1
rlabel polycontact -633 133 -633 133 1 g0
rlabel ndiffusion -651 120 -651 120 1 n31
rlabel ndiffusion -636 120 -636 120 1 n32
rlabel ndcontact -623 119 -623 119 1 nand18
rlabel polycontact -601 136 -601 136 1 nand18
rlabel pdcontact -623 177 -623 177 1 nand18
rlabel pdcontact -652 176 -652 176 1 nand18
rlabel metal1 -587 136 -587 136 1 p2p1g0
rlabel pdcontact -594 155 -594 155 1 p2p1g0
rlabel ndcontact -594 128 -594 128 1 p2p1g0
rlabel polycontact -655 250 -655 250 1 p2
rlabel polycontact -641 242 -641 242 1 g1
rlabel ndiffusion -648 231 -648 231 1 n33
rlabel polycontact -605 242 -605 242 1 nand19
rlabel ndcontact -631 231 -631 231 1 nand19
rlabel pdcontact -648 278 -648 278 1 nand19
rlabel metal1 -592 242 -592 242 1 p2g1
rlabel pdcontact -598 261 -598 261 1 p2g1
rlabel ndcontact -598 234 -598 234 1 p2g1
rlabel polycontact -553 213 -553 213 1 p2g1
rlabel polycontact -529 200 -529 200 1 p2p1g0
rlabel polycontact -542 207 -542 207 1 g2
rlabel metal1 -473 219 -473 219 1 c3
rlabel pdcontact -480 238 -480 238 1 c3
rlabel ndcontact -480 211 -480 211 1 c3
rlabel pdiffusion -545 239 -545 239 1 n34
rlabel pdiffusion -533 238 -533 238 1 n35
rlabel polycontact -487 219 -487 219 1 nor10
rlabel pdcontact -513 239 -513 239 1 nor10
rlabel ndcontact -513 187 -513 187 1 nor10
rlabel polycontact -448 513 -448 513 1 nor11
rlabel pdcontact -474 533 -474 533 1 nor11
rlabel ndcontact -544 187 -544 187 1 nor10
rlabel ndcontact -484 481 -484 481 1 nor11
rlabel ndcontact -505 481 -505 481 1 nor11
rlabel metal1 -434 513 -434 513 7 c4
rlabel ndcontact -441 505 -441 505 1 c4
rlabel pdcontact -441 532 -441 532 1 c4
rlabel ndiffusion -636 355 -636 355 1 n36
rlabel ndiffusion -621 355 -621 355 1 n37
rlabel ndiffusion -614 354 -614 354 1 n38
rlabel ndiffusion -633 477 -633 477 1 n39
rlabel ndiffusion -618 477 -618 477 1 n40
rlabel ndiffusion -630 588 -630 588 1 n41
rlabel pdiffusion -506 533 -506 533 1 n42
rlabel pdiffusion -494 532 -494 532 1 n43
rlabel pdiffusion -484 533 -484 533 1 n44
rlabel polycontact -586 371 -586 371 1 nand20
rlabel ndcontact -603 351 -603 351 1 nand20
rlabel pdcontact -614 412 -614 412 1 nand20
rlabel pdcontact -637 411 -637 411 1 nand20
rlabel ndcontact -605 476 -605 476 1 nand21
rlabel pdcontact -605 534 -605 534 1 nand21
rlabel pdcontact -634 533 -634 533 1 nand21
rlabel polycontact -583 493 -583 493 1 nand21
rlabel polycontact -587 599 -587 599 1 nand22
rlabel ndcontact -613 588 -613 588 1 nand22
rlabel pdcontact -630 635 -630 635 1 nand22
rlabel polycontact -637 607 -637 607 1 p3
rlabel polycontact -623 599 -623 599 1 g2
rlabel metal1 -573 599 -573 599 1 p3g2
rlabel pdcontact -580 618 -580 618 1 p3g2
rlabel ndcontact -580 591 -580 591 1 p3g2
rlabel polycontact -644 506 -644 506 1 p3
rlabel polycontact -631 498 -631 498 1 p2
rlabel polycontact -615 490 -615 490 1 g1
rlabel metal1 -569 493 -569 493 1 p3p2g1
rlabel ndcontact -576 485 -576 485 1 p3p2g1
rlabel pdcontact -576 512 -576 512 1 p3p2g1
rlabel polycontact -647 384 -647 384 1 p3
rlabel polycontact -634 376 -634 376 1 p2
rlabel polycontact -622 370 -622 370 1 p1
rlabel polycontact -611 365 -611 365 1 g0
rlabel metal1 -572 371 -572 371 1 p3p2p1g0
rlabel ndcontact -579 363 -579 363 1 p3p2p1g0
rlabel pdcontact -579 390 -579 390 1 p3p2p1g0
rlabel polycontact -514 507 -514 507 1 p3g2
rlabel polycontact -503 500 -503 500 1 p3p2g1
rlabel polycontact -492 493 -492 493 1 p3p2p1g0
rlabel polycontact -482 494 -482 494 1 g3
rlabel metal1 -290 52 -290 52 5 vdd
rlabel pdcontact -294 39 -294 39 1 vdd
rlabel ndcontact -294 12 -294 12 1 gnd
rlabel metal1 -292 -1 -292 -1 1 gnd
rlabel metal1 -257 53 -257 53 5 vdd
rlabel pdcontact -261 40 -261 40 1 vdd
rlabel ndcontact -261 13 -261 13 1 gnd
rlabel metal1 -259 0 -259 0 1 gnd
rlabel pdcontact -202 40 -202 40 1 vdd
rlabel pdcontact -233 41 -233 41 1 vdd
rlabel ndcontact -233 -3 -233 -3 1 gnd
rlabel metal1 -219 56 -219 56 5 vdd
rlabel metal1 -175 -16 -175 -16 1 gnd
rlabel ndcontact -177 -3 -177 -3 1 gnd
rlabel pdcontact -177 24 -177 24 1 vdd
rlabel pdcontact -116 40 -116 40 1 vdd
rlabel pdcontact -147 41 -147 41 1 vdd
rlabel ndcontact -147 -3 -147 -3 1 gnd
rlabel metal1 -133 56 -133 56 5 vdd
rlabel metal1 -89 -16 -89 -16 1 gnd
rlabel ndcontact -91 -3 -91 -3 1 gnd
rlabel pdcontact -91 24 -91 24 1 vdd
rlabel pdcontact -23 26 -23 26 1 vdd
rlabel ndcontact -23 -1 -23 -1 1 gnd
rlabel metal1 -52 -18 -52 -18 1 gnd
rlabel metal1 -52 47 -52 47 5 vdd
rlabel pdcontact -61 29 -61 29 1 vdd
rlabel ndcontact -43 -8 -43 -8 1 gnd
rlabel ndcontact -61 -7 -61 -7 1 gnd
rlabel metal1 -290 169 -290 169 5 vdd
rlabel pdcontact -294 156 -294 156 1 vdd
rlabel ndcontact -294 129 -294 129 1 gnd
rlabel metal1 -292 116 -292 116 1 gnd
rlabel metal1 -257 170 -257 170 5 vdd
rlabel pdcontact -261 157 -261 157 1 vdd
rlabel ndcontact -261 130 -261 130 1 gnd
rlabel metal1 -259 117 -259 117 1 gnd
rlabel pdcontact -202 157 -202 157 1 vdd
rlabel pdcontact -233 158 -233 158 1 vdd
rlabel ndcontact -233 114 -233 114 1 gnd
rlabel metal1 -219 173 -219 173 5 vdd
rlabel metal1 -175 101 -175 101 1 gnd
rlabel ndcontact -177 114 -177 114 1 gnd
rlabel pdcontact -177 141 -177 141 1 vdd
rlabel pdcontact -116 157 -116 157 1 vdd
rlabel pdcontact -147 158 -147 158 1 vdd
rlabel ndcontact -147 114 -147 114 1 gnd
rlabel metal1 -133 173 -133 173 5 vdd
rlabel metal1 -89 101 -89 101 1 gnd
rlabel ndcontact -91 114 -91 114 1 gnd
rlabel pdcontact -91 141 -91 141 1 vdd
rlabel pdcontact -23 143 -23 143 1 vdd
rlabel ndcontact -23 116 -23 116 1 gnd
rlabel metal1 -52 99 -52 99 1 gnd
rlabel metal1 -52 164 -52 164 5 vdd
rlabel pdcontact -61 146 -61 146 1 vdd
rlabel ndcontact -43 109 -43 109 1 gnd
rlabel ndcontact -61 110 -61 110 1 gnd
rlabel polycontact -293 20 -293 20 1 p0
rlabel metal1 -279 20 -279 20 1 p01
rlabel pdcontact -286 39 -286 39 1 p01
rlabel ndcontact -286 12 -286 12 1 p01
rlabel polycontact -260 21 -260 21 1 c0
rlabel metal1 -246 21 -246 21 1 c01
rlabel pdcontact -253 40 -253 40 1 c01
rlabel ndcontact -253 13 -253 13 1 c01
rlabel polycontact -226 13 -226 13 1 p0
rlabel polycontact -212 5 -212 5 1 c01
rlabel pdcontact -219 41 -219 41 1 nand9
rlabel ndcontact -202 -6 -202 -6 1 nand9
rlabel polycontact -176 5 -176 5 1 nand9
rlabel ndcontact -169 -3 -169 -3 1 p0c01
rlabel metal1 -162 5 -162 5 1 p0c01
rlabel pdcontact -169 24 -169 24 1 p0c01
rlabel polycontact -140 13 -140 13 1 p01
rlabel polycontact -126 5 -126 5 1 c0
rlabel pdcontact -133 41 -133 41 1 nand10
rlabel ndcontact -116 -6 -116 -6 1 nand10
rlabel polycontact -90 5 -90 5 1 nand10
rlabel pdcontact -83 24 -83 24 1 p01c0
rlabel ndcontact -83 -3 -83 -3 1 p01c0
rlabel metal1 -76 5 -76 5 1 p01c0
rlabel polycontact -60 8 -60 8 1 p0c01
rlabel polycontact -49 8 -49 8 1 p01c0
rlabel pdcontact -42 29 -42 29 1 nor5
rlabel ndcontact -52 -8 -52 -8 1 nor5
rlabel polycontact -22 7 -22 7 1 nor5
rlabel pdcontact -15 26 -15 26 1 s0
rlabel metal1 -8 7 -8 7 1 s0
rlabel ndcontact -15 -1 -15 -1 1 s0
rlabel ndiffusion -219 -6 -219 -6 1 n17
rlabel ndiffusion -133 -7 -133 -7 1 n18
rlabel pdiffusion -52 30 -52 30 1 n19
rlabel metal1 -8 124 -8 124 1 s1
rlabel ndcontact -15 116 -15 116 1 s1
rlabel pdcontact -15 143 -15 143 1 s1
rlabel polycontact -22 124 -22 124 1 nor6
rlabel pdcontact -42 146 -42 146 1 nor6
rlabel ndcontact -52 109 -52 109 1 nor6
rlabel polycontact -293 137 -293 137 1 p1
rlabel metal1 -279 137 -279 137 1 p11
rlabel pdcontact -286 156 -286 156 1 p11
rlabel ndcontact -286 129 -286 129 1 p11
rlabel metal1 -246 138 -246 138 1 c11
rlabel ndcontact -253 130 -253 130 1 c11
rlabel pdcontact -253 157 -253 157 1 c11
rlabel pdcontact -219 158 -219 158 1 nand11
rlabel ndcontact -202 111 -202 111 1 nand11
rlabel polycontact -176 122 -176 122 1 nand11
rlabel ndiffusion -219 111 -219 111 1 n20
rlabel ndiffusion -133 110 -133 110 1 n21
rlabel pdiffusion -52 147 -52 147 1 n22
rlabel polycontact -49 125 -49 125 1 p11c1
rlabel polycontact -60 125 -60 125 1 p1c11
rlabel metal1 -76 122 -76 122 1 p11c1
rlabel pdcontact -83 141 -83 141 1 p11c1
rlabel ndcontact -83 114 -83 114 1 p11c1
rlabel polycontact -90 122 -90 122 1 nand12
rlabel pdcontact -133 158 -133 158 1 nand12
rlabel ndcontact -116 111 -116 111 1 nand12
rlabel polycontact -140 130 -140 130 1 p11
rlabel ndcontact -169 114 -169 114 1 p1c11
rlabel metal1 -162 122 -162 122 1 p1c11
rlabel pdcontact -169 141 -169 141 1 p1c11
rlabel polycontact -212 122 -212 122 1 c11
rlabel polycontact -226 130 -226 130 1 p1
rlabel metal1 -288 289 -288 289 5 vdd
rlabel pdcontact -292 276 -292 276 1 vdd
rlabel ndcontact -292 249 -292 249 1 gnd
rlabel metal1 -290 236 -290 236 1 gnd
rlabel metal1 -255 290 -255 290 5 vdd
rlabel pdcontact -259 277 -259 277 1 vdd
rlabel ndcontact -259 250 -259 250 1 gnd
rlabel metal1 -257 237 -257 237 1 gnd
rlabel pdcontact -200 277 -200 277 1 vdd
rlabel pdcontact -231 278 -231 278 1 vdd
rlabel ndcontact -231 234 -231 234 1 gnd
rlabel metal1 -217 293 -217 293 5 vdd
rlabel metal1 -173 221 -173 221 1 gnd
rlabel ndcontact -175 234 -175 234 1 gnd
rlabel pdcontact -175 261 -175 261 1 vdd
rlabel pdcontact -114 277 -114 277 1 vdd
rlabel pdcontact -145 278 -145 278 1 vdd
rlabel ndcontact -145 234 -145 234 1 gnd
rlabel metal1 -131 293 -131 293 5 vdd
rlabel metal1 -87 221 -87 221 1 gnd
rlabel ndcontact -89 234 -89 234 1 gnd
rlabel pdcontact -89 261 -89 261 1 vdd
rlabel pdcontact -21 263 -21 263 1 vdd
rlabel ndcontact -21 236 -21 236 1 gnd
rlabel metal1 -50 219 -50 219 1 gnd
rlabel metal1 -50 284 -50 284 5 vdd
rlabel pdcontact -59 266 -59 266 1 vdd
rlabel ndcontact -41 229 -41 229 1 gnd
rlabel ndcontact -59 230 -59 230 1 gnd
rlabel metal1 -288 406 -288 406 5 vdd
rlabel pdcontact -292 393 -292 393 1 vdd
rlabel ndcontact -292 366 -292 366 1 gnd
rlabel metal1 -290 353 -290 353 1 gnd
rlabel metal1 -255 407 -255 407 5 vdd
rlabel pdcontact -259 394 -259 394 1 vdd
rlabel ndcontact -259 367 -259 367 1 gnd
rlabel metal1 -257 354 -257 354 1 gnd
rlabel pdcontact -200 394 -200 394 1 vdd
rlabel pdcontact -231 395 -231 395 1 vdd
rlabel ndcontact -231 351 -231 351 1 gnd
rlabel metal1 -217 410 -217 410 5 vdd
rlabel metal1 -173 338 -173 338 1 gnd
rlabel ndcontact -175 351 -175 351 1 gnd
rlabel pdcontact -175 378 -175 378 1 vdd
rlabel pdcontact -114 394 -114 394 1 vdd
rlabel pdcontact -145 395 -145 395 1 vdd
rlabel ndcontact -145 351 -145 351 1 gnd
rlabel metal1 -131 410 -131 410 5 vdd
rlabel metal1 -87 338 -87 338 1 gnd
rlabel ndcontact -89 351 -89 351 1 gnd
rlabel pdcontact -89 378 -89 378 1 vdd
rlabel pdcontact -21 380 -21 380 1 vdd
rlabel ndcontact -21 353 -21 353 1 gnd
rlabel metal1 -50 336 -50 336 1 gnd
rlabel metal1 -50 401 -50 401 5 vdd
rlabel pdcontact -59 383 -59 383 1 vdd
rlabel ndcontact -41 346 -41 346 1 gnd
rlabel ndcontact -59 347 -59 347 1 gnd
rlabel metal1 -6 244 -6 244 7 s2
rlabel ndcontact -13 236 -13 236 1 s2
rlabel pdcontact -13 263 -13 263 1 s2
rlabel polycontact -20 244 -20 244 1 nor7
rlabel pdcontact -40 266 -40 266 1 nor7
rlabel ndcontact -50 229 -50 229 1 nor7
rlabel polycontact -47 245 -47 245 1 p21c2
rlabel polycontact -58 245 -58 245 1 p2c21
rlabel ndiffusion -217 231 -217 231 1 n23
rlabel ndiffusion -131 230 -131 230 1 n24
rlabel pdiffusion -50 267 -50 267 1 n25
rlabel metal1 -74 242 -74 242 1 p21c2
rlabel pdcontact -217 278 -217 278 1 nand13
rlabel ndcontact -200 231 -200 231 1 nand13
rlabel polycontact -174 242 -174 242 1 nand13
rlabel polycontact -88 242 -88 242 1 nand14
rlabel ndcontact -114 231 -114 231 1 nand14
rlabel pdcontact -131 278 -131 278 1 nand14
rlabel ndcontact -81 234 -81 234 1 p21c2
rlabel pdcontact -81 261 -81 261 1 p21c2
rlabel polycontact -124 242 -124 242 1 c2
rlabel polycontact -138 250 -138 250 1 p21
rlabel metal1 -160 242 -160 242 1 p2c21
rlabel pdcontact -167 261 -167 261 1 p2c21
rlabel ndcontact -167 234 -167 234 1 p2c21
rlabel polycontact -210 242 -210 242 1 c21
rlabel polycontact -224 250 -224 250 1 p2
rlabel ndcontact -251 250 -251 250 1 c21
rlabel metal1 -244 258 -244 258 1 c21
rlabel pdcontact -251 277 -251 277 1 c21
rlabel polycontact -258 258 -258 258 1 c2
rlabel metal1 -277 257 -277 257 1 p21
rlabel polycontact -291 257 -291 257 1 p2
rlabel pdcontact -284 276 -284 276 1 p21
rlabel ndcontact -284 249 -284 249 1 p21
rlabel polycontact -20 361 -20 361 1 nor8
rlabel ndcontact -50 346 -50 346 1 nor8
rlabel pdcontact -40 383 -40 383 1 nor8
rlabel pdiffusion -50 384 -50 384 1 n26
rlabel ndiffusion -131 347 -131 347 1 n27
rlabel ndiffusion -217 348 -217 348 1 n28
rlabel ndcontact -200 348 -200 348 1 nand15
rlabel polycontact -174 359 -174 359 1 nand15
rlabel pdcontact -217 395 -217 395 1 nand15
rlabel ndcontact -114 348 -114 348 1 nand16
rlabel polycontact -88 359 -88 359 1 nand16
rlabel pdcontact -131 395 -131 395 1 nand16
rlabel metal1 -6 361 -6 361 7 s3
rlabel ndcontact -13 353 -13 353 1 s3
rlabel pdcontact -13 380 -13 380 1 s3
rlabel polycontact -291 374 -291 374 1 p3
rlabel metal1 -277 374 -277 374 1 p31
rlabel polycontact -258 375 -258 375 1 c3
rlabel ndcontact -284 366 -284 366 1 p31
rlabel pdcontact -284 393 -284 393 1 p31
rlabel metal1 -244 375 -244 375 1 c31
rlabel ndcontact -251 367 -251 367 1 c31
rlabel pdcontact -251 394 -251 394 1 c31
rlabel polycontact -224 367 -224 367 1 p3
rlabel polycontact -210 359 -210 359 1 c31
rlabel metal1 -160 359 -160 359 1 p3c31
rlabel ndcontact -167 351 -167 351 1 p3c31
rlabel pdcontact -167 378 -167 378 1 p3c31
rlabel polycontact -138 367 -138 367 1 p31
rlabel polycontact -124 359 -124 359 1 c3
rlabel metal1 -74 359 -74 359 1 p31c3
rlabel ndcontact -81 351 -81 351 1 p31c3
rlabel pdcontact -81 378 -81 378 1 p31c3
rlabel polycontact -58 362 -58 362 1 p3c31
rlabel polycontact -47 362 -47 362 1 p31c3
rlabel polycontact -260 138 -260 138 1 g0
rlabel polycontact -126 122 -126 122 1 g0
rlabel pdcontact -931 33 -931 33 1 vdd
rlabel ndcontact -931 6 -931 6 1 gnd
rlabel metal1 -929 -7 -929 -7 1 gnd
rlabel metal1 -973 65 -973 65 5 vdd
rlabel ndcontact -987 6 -987 6 1 gnd
rlabel pdcontact -987 50 -987 50 1 vdd
rlabel pdcontact -956 49 -956 49 1 vdd
rlabel polycontact -980 22 -980 22 1 a0
rlabel polycontact -966 14 -966 14 1 b0
rlabel pdcontact -973 50 -973 50 1 a0b0
rlabel ndcontact -956 3 -956 3 1 a0b0
rlabel polycontact -930 14 -930 14 1 a0b0
rlabel ndcontact -923 6 -923 6 1 g0
rlabel metal1 -916 14 -916 14 7 g0
rlabel pdcontact -923 33 -923 33 1 g0
rlabel metal1 -1176 149 -1176 149 5 vdd
rlabel pdcontact -1180 136 -1180 136 1 vdd
rlabel ndcontact -1180 109 -1180 109 1 gnd
rlabel metal1 -1178 96 -1178 96 1 gnd
rlabel metal1 -1143 150 -1143 150 5 vdd
rlabel pdcontact -1147 137 -1147 137 1 vdd
rlabel ndcontact -1147 110 -1147 110 1 gnd
rlabel metal1 -1145 97 -1145 97 1 gnd
rlabel ndiffusion -1105 91 -1105 91 1 n1
rlabel pdcontact -1088 137 -1088 137 1 vdd
rlabel pdcontact -1119 138 -1119 138 1 vdd
rlabel ndcontact -1119 94 -1119 94 1 gnd
rlabel metal1 -1105 153 -1105 153 5 vdd
rlabel metal1 -1061 81 -1061 81 1 gnd
rlabel ndcontact -1063 94 -1063 94 1 gnd
rlabel pdcontact -1063 121 -1063 121 1 vdd
rlabel pdcontact -1002 137 -1002 137 1 vdd
rlabel pdcontact -1033 138 -1033 138 1 vdd
rlabel ndcontact -1033 94 -1033 94 1 gnd
rlabel metal1 -1019 153 -1019 153 5 vdd
rlabel metal1 -975 81 -975 81 1 gnd
rlabel ndcontact -977 94 -977 94 1 gnd
rlabel pdcontact -977 121 -977 121 1 vdd
rlabel polycontact -1062 102 -1062 102 1 nand1
rlabel pdcontact -1105 138 -1105 138 1 nand1
rlabel ndiffusion -1019 90 -1019 90 1 n2
rlabel ndcontact -1088 91 -1088 91 1 nand1
rlabel ndcontact -1002 91 -1002 91 1 nand2
rlabel pdcontact -1019 138 -1019 138 1 nand2
rlabel polycontact -976 102 -976 102 1 nand2
rlabel pdcontact -909 123 -909 123 1 vdd
rlabel ndcontact -909 96 -909 96 1 gnd
rlabel metal1 -938 79 -938 79 1 gnd
rlabel metal1 -938 144 -938 144 5 vdd
rlabel pdcontact -947 126 -947 126 1 vdd
rlabel ndcontact -929 89 -929 89 1 gnd
rlabel ndcontact -947 90 -947 90 1 gnd
rlabel pdiffusion -938 127 -938 127 1 n3
rlabel pdcontact -928 126 -928 126 1 nor
rlabel ndcontact -938 89 -938 89 1 nor
rlabel polycontact -908 104 -908 104 1 nor
rlabel polycontact -1179 117 -1179 117 1 a0
rlabel pdcontact -1172 136 -1172 136 1 a01
rlabel metal1 -1165 117 -1165 117 1 a01
rlabel ndcontact -1172 109 -1172 109 1 a01
rlabel polycontact -1146 118 -1146 118 1 b0
rlabel ndcontact -1139 110 -1139 110 1 b01
rlabel metal1 -1132 118 -1132 118 1 b01
rlabel pdcontact -1139 137 -1139 137 1 b01
rlabel polycontact -1112 110 -1112 110 1 a0
rlabel polycontact -1098 102 -1098 102 1 b01
rlabel pdcontact -1055 121 -1055 121 1 a0b01
rlabel metal1 -1048 102 -1048 102 1 a0b01
rlabel ndcontact -1055 94 -1055 94 1 a0b01
rlabel polycontact -1026 110 -1026 110 1 a01
rlabel polycontact -1012 102 -1012 102 1 b0
rlabel pdcontact -969 121 -969 121 1 a01b0
rlabel metal1 -962 102 -962 102 1 a01b0
rlabel ndcontact -969 94 -969 94 1 a01b0
rlabel polycontact -946 105 -946 105 1 a0b01
rlabel polycontact -935 105 -935 105 1 a01b0
rlabel ndiffusion -973 3 -973 3 1 n4
rlabel ndcontact -901 96 -901 96 1 p0
rlabel metal1 -894 104 -894 104 7 p0
rlabel pdcontact -901 123 -901 123 1 p0
rlabel pdcontact -934 261 -934 261 1 vdd
rlabel ndcontact -934 234 -934 234 1 gnd
rlabel metal1 -932 221 -932 221 1 gnd
rlabel metal1 -976 293 -976 293 5 vdd
rlabel ndcontact -990 234 -990 234 1 gnd
rlabel pdcontact -990 278 -990 278 1 vdd
rlabel pdcontact -959 277 -959 277 1 vdd
rlabel metal1 -1179 377 -1179 377 5 vdd
rlabel pdcontact -1183 364 -1183 364 1 vdd
rlabel ndcontact -1183 337 -1183 337 1 gnd
rlabel metal1 -1181 324 -1181 324 1 gnd
rlabel metal1 -1146 378 -1146 378 5 vdd
rlabel pdcontact -1150 365 -1150 365 1 vdd
rlabel ndcontact -1150 338 -1150 338 1 gnd
rlabel metal1 -1148 325 -1148 325 1 gnd
rlabel pdcontact -1091 365 -1091 365 1 vdd
rlabel pdcontact -1122 366 -1122 366 1 vdd
rlabel ndcontact -1122 322 -1122 322 1 gnd
rlabel metal1 -1108 381 -1108 381 5 vdd
rlabel metal1 -1064 309 -1064 309 1 gnd
rlabel ndcontact -1066 322 -1066 322 1 gnd
rlabel pdcontact -1066 349 -1066 349 1 vdd
rlabel pdcontact -1005 365 -1005 365 1 vdd
rlabel pdcontact -1036 366 -1036 366 1 vdd
rlabel ndcontact -1036 322 -1036 322 1 gnd
rlabel metal1 -1022 381 -1022 381 5 vdd
rlabel metal1 -978 309 -978 309 1 gnd
rlabel ndcontact -980 322 -980 322 1 gnd
rlabel pdcontact -980 349 -980 349 1 vdd
rlabel pdcontact -912 351 -912 351 1 vdd
rlabel ndcontact -912 324 -912 324 1 gnd
rlabel metal1 -941 307 -941 307 1 gnd
rlabel metal1 -941 372 -941 372 5 vdd
rlabel pdcontact -950 354 -950 354 1 vdd
rlabel ndcontact -932 317 -932 317 1 gnd
rlabel ndcontact -950 318 -950 318 1 gnd
rlabel pdcontact -933 476 -933 476 1 vdd
rlabel ndcontact -933 449 -933 449 1 gnd
rlabel metal1 -931 436 -931 436 1 gnd
rlabel metal1 -975 508 -975 508 5 vdd
rlabel ndcontact -989 449 -989 449 1 gnd
rlabel pdcontact -989 493 -989 493 1 vdd
rlabel pdcontact -958 492 -958 492 1 vdd
rlabel metal1 -1178 592 -1178 592 5 vdd
rlabel pdcontact -1182 579 -1182 579 1 vdd
rlabel ndcontact -1182 552 -1182 552 1 gnd
rlabel metal1 -1180 539 -1180 539 1 gnd
rlabel metal1 -1145 593 -1145 593 5 vdd
rlabel pdcontact -1149 580 -1149 580 1 vdd
rlabel ndcontact -1149 553 -1149 553 1 gnd
rlabel metal1 -1147 540 -1147 540 1 gnd
rlabel pdcontact -1090 580 -1090 580 1 vdd
rlabel pdcontact -1121 581 -1121 581 1 vdd
rlabel ndcontact -1121 537 -1121 537 1 gnd
rlabel metal1 -1107 596 -1107 596 5 vdd
rlabel metal1 -1063 524 -1063 524 1 gnd
rlabel ndcontact -1065 537 -1065 537 1 gnd
rlabel pdcontact -1065 564 -1065 564 1 vdd
rlabel pdcontact -1004 580 -1004 580 1 vdd
rlabel pdcontact -1035 581 -1035 581 1 vdd
rlabel ndcontact -1035 537 -1035 537 1 gnd
rlabel metal1 -1021 596 -1021 596 5 vdd
rlabel metal1 -977 524 -977 524 1 gnd
rlabel ndcontact -979 537 -979 537 1 gnd
rlabel pdcontact -979 564 -979 564 1 vdd
rlabel pdcontact -911 566 -911 566 1 vdd
rlabel ndcontact -911 539 -911 539 1 gnd
rlabel metal1 -940 522 -940 522 1 gnd
rlabel metal1 -940 587 -940 587 5 vdd
rlabel pdcontact -949 569 -949 569 1 vdd
rlabel ndcontact -931 532 -931 532 1 gnd
rlabel ndcontact -949 533 -949 533 1 gnd
rlabel pdcontact -931 688 -931 688 1 vdd
rlabel ndcontact -931 661 -931 661 1 gnd
rlabel metal1 -929 648 -929 648 1 gnd
rlabel metal1 -973 720 -973 720 5 vdd
rlabel ndcontact -987 661 -987 661 1 gnd
rlabel pdcontact -987 705 -987 705 1 vdd
rlabel pdcontact -956 704 -956 704 1 vdd
rlabel metal1 -1176 804 -1176 804 5 vdd
rlabel pdcontact -1180 791 -1180 791 1 vdd
rlabel ndcontact -1180 764 -1180 764 1 gnd
rlabel metal1 -1178 751 -1178 751 1 gnd
rlabel metal1 -1143 805 -1143 805 5 vdd
rlabel pdcontact -1147 792 -1147 792 1 vdd
rlabel ndcontact -1147 765 -1147 765 1 gnd
rlabel metal1 -1145 752 -1145 752 1 gnd
rlabel pdcontact -1088 792 -1088 792 1 vdd
rlabel pdcontact -1119 793 -1119 793 1 vdd
rlabel ndcontact -1119 749 -1119 749 1 gnd
rlabel metal1 -1105 808 -1105 808 5 vdd
rlabel metal1 -1061 736 -1061 736 1 gnd
rlabel ndcontact -1063 749 -1063 749 1 gnd
rlabel pdcontact -1063 776 -1063 776 1 vdd
rlabel pdcontact -1002 792 -1002 792 1 vdd
rlabel pdcontact -1033 793 -1033 793 1 vdd
rlabel ndcontact -1033 749 -1033 749 1 gnd
rlabel metal1 -1019 808 -1019 808 5 vdd
rlabel metal1 -975 736 -975 736 1 gnd
rlabel ndcontact -977 749 -977 749 1 gnd
rlabel pdcontact -977 776 -977 776 1 vdd
rlabel pdcontact -909 778 -909 778 1 vdd
rlabel ndcontact -909 751 -909 751 1 gnd
rlabel metal1 -938 734 -938 734 1 gnd
rlabel metal1 -938 799 -938 799 5 vdd
rlabel pdcontact -947 781 -947 781 1 vdd
rlabel ndcontact -929 744 -929 744 1 gnd
rlabel ndcontact -947 745 -947 745 1 gnd
rlabel polycontact -983 250 -983 250 1 a1
rlabel polycontact -969 242 -969 242 1 b1
rlabel pdcontact -976 278 -976 278 1 a1b1
rlabel ndcontact -959 231 -959 231 1 a1b1
rlabel polycontact -933 242 -933 242 1 a1b1
rlabel pdcontact -926 261 -926 261 1 g1
rlabel metal1 -919 242 -919 242 1 g1
rlabel ndcontact -904 324 -904 324 1 p1
rlabel metal1 -897 332 -897 332 1 p1
rlabel pdcontact -904 351 -904 351 1 p1
rlabel polycontact -911 332 -911 332 1 nor2
rlabel pdcontact -931 354 -931 354 1 nor2
rlabel ndcontact -941 317 -941 317 1 nor2
rlabel ndiffusion -976 231 -976 231 1 n5
rlabel pdiffusion -941 355 -941 355 1 n6
rlabel ndiffusion -1022 318 -1022 318 1 n7
rlabel ndiffusion -1108 319 -1108 319 1 n8
rlabel polycontact -1182 345 -1182 345 1 a1
rlabel metal1 -1168 345 -1168 345 1 a11
rlabel ndcontact -1175 337 -1175 337 1 a11
rlabel pdcontact -1175 364 -1175 364 1 a11
rlabel polycontact -1149 346 -1149 346 1 b1
rlabel metal1 -1135 346 -1135 346 1 b11
rlabel pdcontact -1142 365 -1142 365 1 b11
rlabel ndcontact -1142 338 -1142 338 1 b11
rlabel pdcontact -1108 366 -1108 366 1 nand3
rlabel ndcontact -1091 319 -1091 319 1 nand3
rlabel polycontact -1065 330 -1065 330 1 nand3
rlabel polycontact -1115 339 -1115 339 1 a1
rlabel polycontact -1101 330 -1101 330 1 b11
rlabel pdcontact -1058 349 -1058 349 1 a1b11
rlabel metal1 -1051 330 -1051 330 1 a1b11
rlabel ndcontact -1058 322 -1058 322 1 a1b11
rlabel polycontact -1029 338 -1029 338 1 a11
rlabel polycontact -1015 330 -1015 330 1 b1
rlabel pdcontact -1022 366 -1022 366 1 nand4
rlabel ndcontact -1005 319 -1005 319 1 nand4
rlabel polycontact -979 330 -979 330 1 nand4
rlabel ndcontact -972 322 -972 322 1 a11b1
rlabel metal1 -965 330 -965 330 1 a11b1
rlabel pdcontact -972 349 -972 349 1 a11b1
rlabel polycontact -949 333 -949 333 1 a1b11
rlabel polycontact -938 333 -938 333 1 a11b1
rlabel ndcontact -925 449 -925 449 1 g2
rlabel metal1 -918 457 -918 457 1 g2
rlabel pdcontact -925 476 -925 476 1 g2
rlabel polycontact -932 457 -932 457 1 a2b2
rlabel ndcontact -958 446 -958 446 1 a2b2
rlabel pdcontact -975 493 -975 493 1 a2b2
rlabel ndiffusion -975 446 -975 446 1 n9
rlabel polycontact -968 457 -968 457 1 b2
rlabel polycontact -982 465 -982 465 1 a2
rlabel polycontact -910 547 -910 547 1 nor3
rlabel pdiffusion -940 570 -940 570 1 n10
rlabel ndiffusion -1021 533 -1021 533 1 n11
rlabel ndiffusion -1107 534 -1107 534 1 n12
rlabel polycontact -1181 560 -1181 560 1 a2
rlabel metal1 -1167 560 -1167 560 1 a21
rlabel ndcontact -1174 552 -1174 552 1 a21
rlabel pdcontact -1174 579 -1174 579 1 a21
rlabel polycontact -1148 561 -1148 561 1 b2
rlabel pdcontact -1141 580 -1141 580 1 b21
rlabel metal1 -1134 561 -1134 561 1 b21
rlabel ndcontact -1141 553 -1141 553 1 b21
rlabel pdcontact -1107 581 -1107 581 1 nand5
rlabel polycontact -1114 553 -1114 553 1 a2
rlabel polycontact -1100 545 -1100 545 1 b21
rlabel ndcontact -1090 534 -1090 534 1 nand5
rlabel polycontact -1064 545 -1064 545 1 nand5
rlabel pdcontact -1057 564 -1057 564 1 a2b21
rlabel ndcontact -1057 537 -1057 537 1 a2b21
rlabel pdcontact -1021 581 -1021 581 1 nand6
rlabel ndcontact -1004 534 -1004 534 1 nand6
rlabel polycontact -1028 553 -1028 553 1 a21
rlabel polycontact -1014 545 -1014 545 1 b2
rlabel polycontact -978 545 -978 545 1 nand6
rlabel ndcontact -971 537 -971 537 1 a21b2
rlabel metal1 -964 545 -964 545 1 a21b2
rlabel pdcontact -971 564 -971 564 1 a21b2
rlabel metal1 -1050 545 -1050 545 1 a2b21
rlabel polycontact -948 548 -948 548 1 a2b21
rlabel polycontact -937 548 -937 548 1 a21b2
rlabel ndcontact -940 532 -940 532 1 nor3
rlabel pdcontact -930 569 -930 569 1 nor3
rlabel polycontact -980 677 -980 677 1 a3
rlabel polycontact -966 669 -966 669 1 b3
rlabel ndiffusion -973 658 -973 658 1 n13
rlabel pdcontact -973 705 -973 705 1 a3b3
rlabel ndcontact -956 658 -956 658 1 a3b3
rlabel polycontact -930 669 -930 669 1 a3b3
rlabel ndcontact -923 661 -923 661 1 g3
rlabel pdcontact -923 688 -923 688 1 g3
rlabel metal1 -916 669 -916 669 1 g3
rlabel metal1 -894 759 -894 759 7 p3
rlabel ndcontact -901 751 -901 751 1 p3
rlabel pdcontact -901 778 -901 778 1 p3
rlabel polycontact -908 759 -908 759 1 nor4
rlabel ndcontact -938 744 -938 744 1 nor4
rlabel pdcontact -928 781 -928 781 1 nor4
rlabel polycontact -935 760 -935 760 1 a31b3
rlabel polycontact -946 760 -946 760 1 a3b31
rlabel pdiffusion -938 782 -938 782 1 n14
rlabel ndcontact -969 749 -969 749 1 a31b3
rlabel metal1 -962 757 -962 757 1 a31b3
rlabel pdcontact -969 776 -969 776 1 a31b3
rlabel ndiffusion -1019 745 -1019 745 1 n15
rlabel ndiffusion -1105 746 -1105 746 1 n16
rlabel polycontact -976 757 -976 757 1 nand7
rlabel ndcontact -1002 746 -1002 746 1 nand7
rlabel pdcontact -1019 793 -1019 793 1 nand7
rlabel polycontact -1062 757 -1062 757 1 nand8
rlabel ndcontact -1088 746 -1088 746 1 nand8
rlabel pdcontact -1105 793 -1105 793 1 nand8
rlabel polycontact -1012 757 -1012 757 1 b3
rlabel polycontact -1026 765 -1026 765 1 a31
rlabel metal1 -1048 757 -1048 757 1 a3b31
rlabel pdcontact -1055 776 -1055 776 1 a3b31
rlabel ndcontact -1055 749 -1055 749 1 a3b31
rlabel polycontact -1112 765 -1112 765 1 a3
rlabel polycontact -1098 757 -1098 757 1 b31
rlabel metal1 -1132 773 -1132 773 1 b31
rlabel polycontact -1146 773 -1146 773 1 b3
rlabel pdcontact -1139 792 -1139 792 1 b31
rlabel ndcontact -1139 765 -1139 765 1 b31
rlabel polycontact -1179 772 -1179 772 1 a3
rlabel metal1 -1165 772 -1165 772 1 a31
rlabel ndcontact -1172 764 -1172 764 1 a31
rlabel pdcontact -1172 791 -1172 791 1 a31
rlabel ndcontact -926 234 -926 234 1 g1
rlabel ndcontact -903 539 -903 539 1 p2
rlabel metal1 -896 547 -896 547 1 p2
rlabel pdcontact -903 566 -903 566 1 p2
<< end >>
