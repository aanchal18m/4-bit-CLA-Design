magic
tech scmos
timestamp 1732085619
<< nwell >>
rect -2164 804 -2054 836
rect -2047 806 -2023 832
rect -1846 794 -1794 797
rect -1905 767 -1881 793
rect -1872 768 -1794 794
rect -1760 778 -1708 797
rect -1672 780 -1637 788
rect -1846 762 -1794 768
rect -1788 762 -1708 778
rect -1788 752 -1764 762
rect -1702 752 -1678 778
rect -1672 755 -1610 780
rect -1634 754 -1610 755
rect -2162 703 -2052 735
rect -2045 705 -2021 731
rect -1714 674 -1662 709
rect -1656 664 -1632 690
rect -2175 578 -2065 610
rect -2058 580 -2034 606
rect -1371 604 -1319 639
rect -1313 594 -1289 620
rect -1848 582 -1796 585
rect -1907 555 -1883 581
rect -1874 556 -1796 582
rect -1762 566 -1710 585
rect -1674 568 -1639 576
rect -1848 550 -1796 556
rect -1790 550 -1710 566
rect -1790 540 -1766 550
rect -1704 540 -1680 566
rect -1674 543 -1612 568
rect -1636 542 -1612 543
rect -1375 518 -1313 538
rect -1240 534 -1179 554
rect -1375 514 -1288 518
rect -1375 503 -1285 514
rect -2175 439 -2065 471
rect -2058 441 -2034 467
rect -1716 462 -1664 497
rect -1309 488 -1285 503
rect -1240 508 -1150 534
rect -1240 502 -1179 508
rect -1658 452 -1634 478
rect -550 456 -440 488
rect -433 458 -409 484
rect -1378 396 -1313 416
rect -958 396 -906 399
rect -1378 392 -1291 396
rect -1378 381 -1288 392
rect -1849 367 -1797 370
rect -2183 331 -2073 363
rect -2066 333 -2042 359
rect -1908 340 -1884 366
rect -1875 341 -1797 367
rect -1763 351 -1711 370
rect -1312 366 -1288 381
rect -1017 369 -993 395
rect -984 370 -906 396
rect -872 380 -820 399
rect -784 382 -749 390
rect -958 364 -906 370
rect -900 364 -820 380
rect -1675 353 -1640 361
rect -900 354 -876 364
rect -814 354 -790 380
rect -784 357 -722 382
rect -746 356 -722 357
rect -548 355 -438 387
rect -431 357 -407 383
rect -1849 335 -1797 341
rect -1791 335 -1711 351
rect -1791 325 -1767 335
rect -1705 325 -1681 351
rect -1675 328 -1613 353
rect -1637 327 -1613 328
rect -2189 222 -2079 254
rect -2072 224 -2048 250
rect -1717 247 -1665 282
rect -1659 237 -1635 263
rect -1389 247 -1337 282
rect -958 279 -906 282
rect -1331 237 -1307 263
rect -1279 240 -1218 253
rect -1017 252 -993 278
rect -984 253 -906 279
rect -872 263 -820 282
rect -784 265 -749 273
rect -958 247 -906 253
rect -900 247 -820 263
rect -1279 214 -1189 240
rect -900 237 -876 247
rect -814 237 -790 263
rect -784 240 -722 265
rect -746 239 -722 240
rect -561 230 -451 262
rect -444 232 -420 258
rect -1279 208 -1218 214
rect -1393 161 -1331 181
rect -1393 157 -1306 161
rect -960 159 -908 162
rect -1393 146 -1303 157
rect -1846 139 -1794 142
rect -2183 94 -2073 126
rect -2066 96 -2042 122
rect -1905 112 -1881 138
rect -1872 113 -1794 139
rect -1760 123 -1708 142
rect -1672 125 -1637 133
rect -1327 131 -1303 146
rect -1019 132 -995 158
rect -986 133 -908 159
rect -874 143 -822 162
rect -786 145 -751 153
rect -960 127 -908 133
rect -902 127 -822 143
rect -1846 107 -1794 113
rect -1788 107 -1708 123
rect -1788 97 -1764 107
rect -1702 97 -1678 123
rect -1672 100 -1610 125
rect -902 117 -878 127
rect -816 117 -792 143
rect -786 120 -724 145
rect -748 119 -724 120
rect -1634 99 -1610 100
rect -561 91 -451 123
rect -444 93 -420 119
rect -1714 19 -1662 54
rect -1656 9 -1632 35
rect -1392 26 -1340 61
rect -1297 49 -1262 57
rect -1334 16 -1310 42
rect -1297 24 -1235 49
rect -960 42 -908 45
rect -1259 23 -1235 24
rect -1019 15 -995 41
rect -986 16 -908 42
rect -874 26 -822 45
rect -786 28 -751 36
rect -960 10 -908 16
rect -902 10 -822 26
rect -902 0 -878 10
rect -816 0 -792 26
rect -786 3 -724 28
rect -748 2 -724 3
rect -569 -17 -459 15
rect -452 -15 -428 11
rect -2187 -52 -2077 -20
rect -2070 -50 -2046 -24
rect -2160 -180 -2050 -148
rect -2043 -178 -2019 -152
<< ntransistor >>
rect -2036 792 -2034 797
rect -2153 786 -2151 791
rect -2121 781 -2119 791
rect -2110 781 -2108 791
rect -2084 781 -2082 791
rect -2073 781 -2071 791
rect -1894 753 -1892 758
rect -1861 754 -1859 759
rect -1830 732 -1827 742
rect -1816 732 -1813 742
rect -1777 738 -1775 743
rect -1744 732 -1741 742
rect -1730 732 -1727 742
rect -1691 738 -1689 743
rect -1623 740 -1621 745
rect -1661 733 -1659 738
rect -1650 733 -1648 738
rect -2034 691 -2032 696
rect -2151 685 -2149 690
rect -2119 680 -2117 690
rect -2108 680 -2106 690
rect -2082 680 -2080 690
rect -2071 680 -2069 690
rect -1698 644 -1695 654
rect -1684 644 -1681 654
rect -1645 650 -1643 655
rect -2047 566 -2045 571
rect -2164 560 -2162 565
rect -2132 555 -2130 565
rect -2121 555 -2119 565
rect -2095 555 -2093 565
rect -2084 555 -2082 565
rect -1355 574 -1352 584
rect -1341 574 -1338 584
rect -1302 580 -1300 585
rect -1896 541 -1894 546
rect -1863 542 -1861 547
rect -1832 520 -1829 530
rect -1818 520 -1815 530
rect -1779 526 -1777 531
rect -1746 520 -1743 530
rect -1732 520 -1729 530
rect -1693 526 -1691 531
rect -1625 528 -1623 533
rect -1663 521 -1661 526
rect -1652 521 -1650 526
rect -1359 460 -1356 475
rect -1345 460 -1342 475
rect -1330 460 -1327 475
rect -1298 474 -1296 479
rect -1163 494 -1161 499
rect -1229 468 -1227 473
rect -1218 468 -1216 473
rect -1207 468 -1205 473
rect -1197 468 -1195 473
rect -422 444 -420 449
rect -1700 432 -1697 442
rect -1686 432 -1683 442
rect -1647 438 -1645 443
rect -539 438 -537 443
rect -507 433 -505 443
rect -496 433 -494 443
rect -470 433 -468 443
rect -459 433 -457 443
rect -2047 427 -2045 432
rect -2164 421 -2162 426
rect -2132 416 -2130 426
rect -2121 416 -2119 426
rect -2095 416 -2093 426
rect -2084 416 -2082 426
rect -1897 326 -1895 331
rect -1864 327 -1862 332
rect -2055 319 -2053 324
rect -2172 313 -2170 318
rect -2140 308 -2138 318
rect -2129 308 -2127 318
rect -2103 308 -2101 318
rect -2092 308 -2090 318
rect -1833 305 -1830 315
rect -1819 305 -1816 315
rect -1780 311 -1778 316
rect -1747 305 -1744 315
rect -1733 305 -1730 315
rect -1694 311 -1692 316
rect -1362 333 -1359 353
rect -1348 333 -1345 353
rect -1337 333 -1334 353
rect -1328 333 -1325 353
rect -1301 352 -1299 357
rect -1006 355 -1004 360
rect -973 356 -971 361
rect -942 334 -939 344
rect -928 334 -925 344
rect -889 340 -887 345
rect -856 334 -853 344
rect -842 334 -839 344
rect -803 340 -801 345
rect -735 342 -733 347
rect -420 343 -418 348
rect -773 335 -771 340
rect -762 335 -760 340
rect -537 337 -535 342
rect -505 332 -503 342
rect -494 332 -492 342
rect -468 332 -466 342
rect -457 332 -455 342
rect -1626 313 -1624 318
rect -1664 306 -1662 311
rect -1653 306 -1651 311
rect -1701 217 -1698 227
rect -1687 217 -1684 227
rect -1648 223 -1646 228
rect -1373 217 -1370 227
rect -1359 217 -1356 227
rect -1320 223 -1318 228
rect -2061 210 -2059 215
rect -1006 238 -1004 243
rect -973 239 -971 244
rect -2178 204 -2176 209
rect -2146 199 -2144 209
rect -2135 199 -2133 209
rect -2109 199 -2107 209
rect -2098 199 -2096 209
rect -942 217 -939 227
rect -928 217 -925 227
rect -889 223 -887 228
rect -856 217 -853 227
rect -842 217 -839 227
rect -803 223 -801 228
rect -735 225 -733 230
rect -773 218 -771 223
rect -762 218 -760 223
rect -433 218 -431 223
rect -550 212 -548 217
rect -518 207 -516 217
rect -507 207 -505 217
rect -481 207 -479 217
rect -470 207 -468 217
rect -1202 200 -1200 205
rect -1268 176 -1266 180
rect -1257 176 -1255 180
rect -1244 176 -1242 180
rect -1894 98 -1892 103
rect -1861 99 -1859 104
rect -2055 82 -2053 87
rect -2172 76 -2170 81
rect -2140 71 -2138 81
rect -2129 71 -2127 81
rect -2103 71 -2101 81
rect -2092 71 -2090 81
rect -1830 77 -1827 87
rect -1816 77 -1813 87
rect -1777 83 -1775 88
rect -1744 77 -1741 87
rect -1730 77 -1727 87
rect -1691 83 -1689 88
rect -1377 103 -1374 118
rect -1363 103 -1360 118
rect -1348 103 -1345 118
rect -1316 117 -1314 122
rect -1008 118 -1006 123
rect -975 119 -973 124
rect -944 97 -941 107
rect -930 97 -927 107
rect -891 103 -889 108
rect -858 97 -855 107
rect -844 97 -841 107
rect -805 103 -803 108
rect -737 105 -735 110
rect -775 98 -773 103
rect -764 98 -762 103
rect -1623 85 -1621 90
rect -1661 78 -1659 83
rect -1650 78 -1648 83
rect -433 79 -431 84
rect -550 73 -548 78
rect -518 68 -516 78
rect -507 68 -505 78
rect -481 68 -479 78
rect -470 68 -468 78
rect -1248 9 -1246 14
rect -1698 -11 -1695 -1
rect -1684 -11 -1681 -1
rect -1645 -5 -1643 0
rect -1376 -4 -1373 6
rect -1362 -4 -1359 6
rect -1323 2 -1321 7
rect -1286 2 -1284 7
rect -1275 2 -1273 7
rect -1008 1 -1006 6
rect -975 2 -973 7
rect -944 -20 -941 -10
rect -930 -20 -927 -10
rect -891 -14 -889 -9
rect -858 -20 -855 -10
rect -844 -20 -841 -10
rect -805 -14 -803 -9
rect -737 -12 -735 -7
rect -775 -19 -773 -14
rect -764 -19 -762 -14
rect -441 -29 -439 -24
rect -558 -35 -556 -30
rect -526 -40 -524 -30
rect -515 -40 -513 -30
rect -489 -40 -487 -30
rect -478 -40 -476 -30
rect -2059 -64 -2057 -59
rect -2176 -70 -2174 -65
rect -2144 -75 -2142 -65
rect -2133 -75 -2131 -65
rect -2107 -75 -2105 -65
rect -2096 -75 -2094 -65
rect -2032 -192 -2030 -187
rect -2149 -198 -2147 -193
rect -2117 -203 -2115 -193
rect -2106 -203 -2104 -193
rect -2080 -203 -2078 -193
rect -2069 -203 -2067 -193
<< ptransistor >>
rect -2153 810 -2151 830
rect -2143 810 -2141 830
rect -2121 815 -2119 825
rect -2084 815 -2082 825
rect -2036 816 -2034 826
rect -1894 777 -1892 787
rect -1861 778 -1859 788
rect -1830 779 -1827 789
rect -1816 779 -1813 789
rect -1744 779 -1741 789
rect -1730 779 -1727 789
rect -1777 762 -1775 772
rect -1691 762 -1689 772
rect -1661 762 -1659 782
rect -1650 762 -1648 782
rect -1623 764 -1621 774
rect -2151 709 -2149 729
rect -2141 709 -2139 729
rect -2119 714 -2117 724
rect -2082 714 -2080 724
rect -2034 715 -2032 725
rect -1698 691 -1695 701
rect -1684 691 -1681 701
rect -1645 674 -1643 684
rect -1355 621 -1352 631
rect -1341 621 -1338 631
rect -2164 584 -2162 604
rect -2154 584 -2152 604
rect -2132 589 -2130 599
rect -2095 589 -2093 599
rect -2047 590 -2045 600
rect -1302 604 -1300 614
rect -1896 565 -1894 575
rect -1863 566 -1861 576
rect -1832 567 -1829 577
rect -1818 567 -1815 577
rect -1746 567 -1743 577
rect -1732 567 -1729 577
rect -1779 550 -1777 560
rect -1693 550 -1691 560
rect -1663 550 -1661 570
rect -1652 550 -1650 570
rect -1625 552 -1623 562
rect -1359 520 -1356 530
rect -1345 520 -1342 530
rect -1330 520 -1327 530
rect -1700 479 -1697 489
rect -1686 479 -1683 489
rect -2164 445 -2162 465
rect -2154 445 -2152 465
rect -2132 450 -2130 460
rect -2095 450 -2093 460
rect -2047 451 -2045 461
rect -1229 508 -1227 548
rect -1218 508 -1216 548
rect -1207 508 -1205 548
rect -1197 508 -1195 548
rect -1163 518 -1161 528
rect -1298 498 -1296 508
rect -1647 462 -1645 472
rect -539 462 -537 482
rect -529 462 -527 482
rect -507 467 -505 477
rect -470 467 -468 477
rect -422 468 -420 478
rect -1362 398 -1359 408
rect -1348 398 -1345 408
rect -1337 398 -1334 408
rect -1328 398 -1325 408
rect -2172 337 -2170 357
rect -2162 337 -2160 357
rect -2140 342 -2138 352
rect -2103 342 -2101 352
rect -2055 343 -2053 353
rect -1897 350 -1895 360
rect -1864 351 -1862 361
rect -1833 352 -1830 362
rect -1819 352 -1816 362
rect -1747 352 -1744 362
rect -1733 352 -1730 362
rect -1780 335 -1778 345
rect -1694 335 -1692 345
rect -1664 335 -1662 355
rect -1653 335 -1651 355
rect -1301 376 -1299 386
rect -1006 379 -1004 389
rect -973 380 -971 390
rect -942 381 -939 391
rect -928 381 -925 391
rect -856 381 -853 391
rect -842 381 -839 391
rect -1626 337 -1624 347
rect -889 364 -887 374
rect -803 364 -801 374
rect -773 364 -771 384
rect -762 364 -760 384
rect -735 366 -733 376
rect -537 361 -535 381
rect -527 361 -525 381
rect -505 366 -503 376
rect -468 366 -466 376
rect -420 367 -418 377
rect -1701 264 -1698 274
rect -1687 264 -1684 274
rect -1373 264 -1370 274
rect -1359 264 -1356 274
rect -2178 228 -2176 248
rect -2168 228 -2166 248
rect -2146 233 -2144 243
rect -2109 233 -2107 243
rect -2061 234 -2059 244
rect -1648 247 -1646 257
rect -1006 262 -1004 272
rect -973 263 -971 273
rect -942 264 -939 274
rect -928 264 -925 274
rect -856 264 -853 274
rect -842 264 -839 274
rect -1320 247 -1318 257
rect -1268 215 -1266 245
rect -1257 215 -1255 245
rect -1244 215 -1242 245
rect -1202 224 -1200 234
rect -889 247 -887 257
rect -803 247 -801 257
rect -773 247 -771 267
rect -762 247 -760 267
rect -735 249 -733 259
rect -550 236 -548 256
rect -540 236 -538 256
rect -518 241 -516 251
rect -481 241 -479 251
rect -433 242 -431 252
rect -1377 163 -1374 173
rect -1363 163 -1360 173
rect -1348 163 -1345 173
rect -1894 122 -1892 132
rect -1861 123 -1859 133
rect -1830 124 -1827 134
rect -1816 124 -1813 134
rect -1744 124 -1741 134
rect -1730 124 -1727 134
rect -2172 100 -2170 120
rect -2162 100 -2160 120
rect -2140 105 -2138 115
rect -2103 105 -2101 115
rect -2055 106 -2053 116
rect -1777 107 -1775 117
rect -1691 107 -1689 117
rect -1661 107 -1659 127
rect -1650 107 -1648 127
rect -1623 109 -1621 119
rect -1316 141 -1314 151
rect -1008 142 -1006 152
rect -975 143 -973 153
rect -944 144 -941 154
rect -930 144 -927 154
rect -858 144 -855 154
rect -844 144 -841 154
rect -891 127 -889 137
rect -805 127 -803 137
rect -775 127 -773 147
rect -764 127 -762 147
rect -737 129 -735 139
rect -550 97 -548 117
rect -540 97 -538 117
rect -518 102 -516 112
rect -481 102 -479 112
rect -433 103 -431 113
rect -1698 36 -1695 46
rect -1684 36 -1681 46
rect -1376 43 -1373 53
rect -1362 43 -1359 53
rect -1645 19 -1643 29
rect -1323 26 -1321 36
rect -1286 31 -1284 51
rect -1275 31 -1273 51
rect -1248 33 -1246 43
rect -1008 25 -1006 35
rect -975 26 -973 36
rect -944 27 -941 37
rect -930 27 -927 37
rect -858 27 -855 37
rect -844 27 -841 37
rect -891 10 -889 20
rect -805 10 -803 20
rect -775 10 -773 30
rect -764 10 -762 30
rect -737 12 -735 22
rect -558 -11 -556 9
rect -548 -11 -546 9
rect -526 -6 -524 4
rect -489 -6 -487 4
rect -441 -5 -439 5
rect -2176 -46 -2174 -26
rect -2166 -46 -2164 -26
rect -2144 -41 -2142 -31
rect -2107 -41 -2105 -31
rect -2059 -40 -2057 -30
rect -2149 -174 -2147 -154
rect -2139 -174 -2137 -154
rect -2117 -169 -2115 -159
rect -2080 -169 -2078 -159
rect -2032 -168 -2030 -158
<< ndiffusion >>
rect -2037 792 -2036 797
rect -2034 792 -2033 797
rect -2154 786 -2153 791
rect -2151 786 -2138 791
rect -2122 781 -2121 791
rect -2119 781 -2110 791
rect -2108 781 -2103 791
rect -2086 781 -2084 791
rect -2082 781 -2073 791
rect -2071 781 -2067 791
rect -1895 753 -1894 758
rect -1892 753 -1891 758
rect -1862 754 -1861 759
rect -1859 754 -1858 759
rect -1833 732 -1830 742
rect -1827 732 -1816 742
rect -1813 732 -1807 742
rect -1778 738 -1777 743
rect -1775 738 -1774 743
rect -1747 732 -1744 742
rect -1741 732 -1730 742
rect -1727 732 -1721 742
rect -1692 738 -1691 743
rect -1689 738 -1688 743
rect -1624 740 -1623 745
rect -1621 740 -1620 745
rect -1662 733 -1661 738
rect -1659 733 -1657 738
rect -1653 733 -1650 738
rect -1648 733 -1647 738
rect -2035 691 -2034 696
rect -2032 691 -2031 696
rect -2152 685 -2151 690
rect -2149 685 -2136 690
rect -2120 680 -2119 690
rect -2117 680 -2108 690
rect -2106 680 -2101 690
rect -2084 680 -2082 690
rect -2080 680 -2071 690
rect -2069 680 -2065 690
rect -1701 644 -1698 654
rect -1695 644 -1684 654
rect -1681 644 -1675 654
rect -1646 650 -1645 655
rect -1643 650 -1642 655
rect -2048 566 -2047 571
rect -2045 566 -2044 571
rect -2165 560 -2164 565
rect -2162 560 -2149 565
rect -2133 555 -2132 565
rect -2130 555 -2121 565
rect -2119 555 -2114 565
rect -2097 555 -2095 565
rect -2093 555 -2084 565
rect -2082 555 -2078 565
rect -1358 574 -1355 584
rect -1352 574 -1341 584
rect -1338 574 -1332 584
rect -1303 580 -1302 585
rect -1300 580 -1299 585
rect -1897 541 -1896 546
rect -1894 541 -1893 546
rect -1864 542 -1863 547
rect -1861 542 -1860 547
rect -1835 520 -1832 530
rect -1829 520 -1818 530
rect -1815 520 -1809 530
rect -1780 526 -1779 531
rect -1777 526 -1776 531
rect -1749 520 -1746 530
rect -1743 520 -1732 530
rect -1729 520 -1723 530
rect -1694 526 -1693 531
rect -1691 526 -1690 531
rect -1626 528 -1625 533
rect -1623 528 -1622 533
rect -1664 521 -1663 526
rect -1661 521 -1659 526
rect -1655 521 -1652 526
rect -1650 521 -1649 526
rect -1363 460 -1359 475
rect -1356 460 -1345 475
rect -1342 460 -1330 475
rect -1327 460 -1324 475
rect -1299 474 -1298 479
rect -1296 474 -1295 479
rect -1164 494 -1163 499
rect -1161 494 -1160 499
rect -1230 468 -1229 473
rect -1227 468 -1224 473
rect -1220 468 -1218 473
rect -1216 468 -1212 473
rect -1208 468 -1207 473
rect -1205 468 -1203 473
rect -1199 468 -1197 473
rect -1195 468 -1194 473
rect -423 444 -422 449
rect -420 444 -419 449
rect -1703 432 -1700 442
rect -1697 432 -1686 442
rect -1683 432 -1677 442
rect -1648 438 -1647 443
rect -1645 438 -1644 443
rect -540 438 -539 443
rect -537 438 -524 443
rect -508 433 -507 443
rect -505 433 -496 443
rect -494 433 -489 443
rect -472 433 -470 443
rect -468 433 -459 443
rect -457 433 -453 443
rect -2048 427 -2047 432
rect -2045 427 -2044 432
rect -2165 421 -2164 426
rect -2162 421 -2149 426
rect -2133 416 -2132 426
rect -2130 416 -2121 426
rect -2119 416 -2114 426
rect -2097 416 -2095 426
rect -2093 416 -2084 426
rect -2082 416 -2078 426
rect -1898 326 -1897 331
rect -1895 326 -1894 331
rect -1865 327 -1864 332
rect -1862 327 -1861 332
rect -2056 319 -2055 324
rect -2053 319 -2052 324
rect -2173 313 -2172 318
rect -2170 313 -2157 318
rect -2141 308 -2140 318
rect -2138 308 -2129 318
rect -2127 308 -2122 318
rect -2105 308 -2103 318
rect -2101 308 -2092 318
rect -2090 308 -2086 318
rect -1836 305 -1833 315
rect -1830 305 -1819 315
rect -1816 305 -1810 315
rect -1781 311 -1780 316
rect -1778 311 -1777 316
rect -1750 305 -1747 315
rect -1744 305 -1733 315
rect -1730 305 -1724 315
rect -1695 311 -1694 316
rect -1692 311 -1691 316
rect -1366 333 -1362 353
rect -1359 333 -1348 353
rect -1345 333 -1337 353
rect -1334 333 -1328 353
rect -1325 333 -1322 353
rect -1302 352 -1301 357
rect -1299 352 -1298 357
rect -1007 355 -1006 360
rect -1004 355 -1003 360
rect -974 356 -973 361
rect -971 356 -970 361
rect -945 334 -942 344
rect -939 334 -928 344
rect -925 334 -919 344
rect -890 340 -889 345
rect -887 340 -886 345
rect -859 334 -856 344
rect -853 334 -842 344
rect -839 334 -833 344
rect -804 340 -803 345
rect -801 340 -800 345
rect -736 342 -735 347
rect -733 342 -732 347
rect -421 343 -420 348
rect -418 343 -417 348
rect -774 335 -773 340
rect -771 335 -769 340
rect -765 335 -762 340
rect -760 335 -759 340
rect -538 337 -537 342
rect -535 337 -522 342
rect -506 332 -505 342
rect -503 332 -494 342
rect -492 332 -487 342
rect -470 332 -468 342
rect -466 332 -457 342
rect -455 332 -451 342
rect -1627 313 -1626 318
rect -1624 313 -1623 318
rect -1665 306 -1664 311
rect -1662 306 -1660 311
rect -1656 306 -1653 311
rect -1651 306 -1650 311
rect -1704 217 -1701 227
rect -1698 217 -1687 227
rect -1684 217 -1678 227
rect -1649 223 -1648 228
rect -1646 223 -1645 228
rect -1376 217 -1373 227
rect -1370 217 -1359 227
rect -1356 217 -1350 227
rect -1321 223 -1320 228
rect -1318 223 -1317 228
rect -2062 210 -2061 215
rect -2059 210 -2058 215
rect -1007 238 -1006 243
rect -1004 238 -1003 243
rect -974 239 -973 244
rect -971 239 -970 244
rect -2179 204 -2178 209
rect -2176 204 -2163 209
rect -2147 199 -2146 209
rect -2144 199 -2135 209
rect -2133 199 -2128 209
rect -2111 199 -2109 209
rect -2107 199 -2098 209
rect -2096 199 -2092 209
rect -945 217 -942 227
rect -939 217 -928 227
rect -925 217 -919 227
rect -890 223 -889 228
rect -887 223 -886 228
rect -859 217 -856 227
rect -853 217 -842 227
rect -839 217 -833 227
rect -804 223 -803 228
rect -801 223 -800 228
rect -736 225 -735 230
rect -733 225 -732 230
rect -774 218 -773 223
rect -771 218 -769 223
rect -765 218 -762 223
rect -760 218 -759 223
rect -434 218 -433 223
rect -431 218 -430 223
rect -551 212 -550 217
rect -548 212 -535 217
rect -519 207 -518 217
rect -516 207 -507 217
rect -505 207 -500 217
rect -483 207 -481 217
rect -479 207 -470 217
rect -468 207 -464 217
rect -1203 200 -1202 205
rect -1200 200 -1199 205
rect -1269 176 -1268 180
rect -1266 176 -1263 180
rect -1259 176 -1257 180
rect -1255 176 -1251 180
rect -1247 176 -1244 180
rect -1242 176 -1233 180
rect -1895 98 -1894 103
rect -1892 98 -1891 103
rect -1862 99 -1861 104
rect -1859 99 -1858 104
rect -2056 82 -2055 87
rect -2053 82 -2052 87
rect -2173 76 -2172 81
rect -2170 76 -2157 81
rect -2141 71 -2140 81
rect -2138 71 -2129 81
rect -2127 71 -2122 81
rect -2105 71 -2103 81
rect -2101 71 -2092 81
rect -2090 71 -2086 81
rect -1833 77 -1830 87
rect -1827 77 -1816 87
rect -1813 77 -1807 87
rect -1778 83 -1777 88
rect -1775 83 -1774 88
rect -1747 77 -1744 87
rect -1741 77 -1730 87
rect -1727 77 -1721 87
rect -1692 83 -1691 88
rect -1689 83 -1688 88
rect -1381 103 -1377 118
rect -1374 103 -1363 118
rect -1360 103 -1348 118
rect -1345 103 -1342 118
rect -1317 117 -1316 122
rect -1314 117 -1313 122
rect -1009 118 -1008 123
rect -1006 118 -1005 123
rect -976 119 -975 124
rect -973 119 -972 124
rect -947 97 -944 107
rect -941 97 -930 107
rect -927 97 -921 107
rect -892 103 -891 108
rect -889 103 -888 108
rect -861 97 -858 107
rect -855 97 -844 107
rect -841 97 -835 107
rect -806 103 -805 108
rect -803 103 -802 108
rect -738 105 -737 110
rect -735 105 -734 110
rect -776 98 -775 103
rect -773 98 -771 103
rect -767 98 -764 103
rect -762 98 -761 103
rect -1624 85 -1623 90
rect -1621 85 -1620 90
rect -1662 78 -1661 83
rect -1659 78 -1657 83
rect -1653 78 -1650 83
rect -1648 78 -1647 83
rect -434 79 -433 84
rect -431 79 -430 84
rect -551 73 -550 78
rect -548 73 -535 78
rect -519 68 -518 78
rect -516 68 -507 78
rect -505 68 -500 78
rect -483 68 -481 78
rect -479 68 -470 78
rect -468 68 -464 78
rect -1249 9 -1248 14
rect -1246 9 -1245 14
rect -1701 -11 -1698 -1
rect -1695 -11 -1684 -1
rect -1681 -11 -1675 -1
rect -1646 -5 -1645 0
rect -1643 -5 -1642 0
rect -1379 -4 -1376 6
rect -1373 -4 -1362 6
rect -1359 -4 -1353 6
rect -1324 2 -1323 7
rect -1321 2 -1320 7
rect -1287 2 -1286 7
rect -1284 2 -1282 7
rect -1278 2 -1275 7
rect -1273 2 -1272 7
rect -1009 1 -1008 6
rect -1006 1 -1005 6
rect -976 2 -975 7
rect -973 2 -972 7
rect -947 -20 -944 -10
rect -941 -20 -930 -10
rect -927 -20 -921 -10
rect -892 -14 -891 -9
rect -889 -14 -888 -9
rect -861 -20 -858 -10
rect -855 -20 -844 -10
rect -841 -20 -835 -10
rect -806 -14 -805 -9
rect -803 -14 -802 -9
rect -738 -12 -737 -7
rect -735 -12 -734 -7
rect -776 -19 -775 -14
rect -773 -19 -771 -14
rect -767 -19 -764 -14
rect -762 -19 -761 -14
rect -442 -29 -441 -24
rect -439 -29 -438 -24
rect -559 -35 -558 -30
rect -556 -35 -543 -30
rect -527 -40 -526 -30
rect -524 -40 -515 -30
rect -513 -40 -508 -30
rect -491 -40 -489 -30
rect -487 -40 -478 -30
rect -476 -40 -472 -30
rect -2060 -64 -2059 -59
rect -2057 -64 -2056 -59
rect -2177 -70 -2176 -65
rect -2174 -70 -2161 -65
rect -2145 -75 -2144 -65
rect -2142 -75 -2133 -65
rect -2131 -75 -2126 -65
rect -2109 -75 -2107 -65
rect -2105 -75 -2096 -65
rect -2094 -75 -2090 -65
rect -2033 -192 -2032 -187
rect -2030 -192 -2029 -187
rect -2150 -198 -2149 -193
rect -2147 -198 -2134 -193
rect -2118 -203 -2117 -193
rect -2115 -203 -2106 -193
rect -2104 -203 -2099 -193
rect -2082 -203 -2080 -193
rect -2078 -203 -2069 -193
rect -2067 -203 -2063 -193
<< pdiffusion >>
rect -2154 810 -2153 830
rect -2151 810 -2143 830
rect -2141 810 -2138 830
rect -2122 815 -2121 825
rect -2119 815 -2103 825
rect -2086 815 -2084 825
rect -2082 815 -2067 825
rect -2037 816 -2036 826
rect -2034 816 -2033 826
rect -1895 777 -1894 787
rect -1892 777 -1891 787
rect -1862 778 -1861 788
rect -1859 778 -1858 788
rect -1833 779 -1830 789
rect -1827 779 -1824 789
rect -1819 779 -1816 789
rect -1813 779 -1807 789
rect -1747 779 -1744 789
rect -1741 779 -1738 789
rect -1733 779 -1730 789
rect -1727 779 -1721 789
rect -1778 762 -1777 772
rect -1775 762 -1774 772
rect -1692 762 -1691 772
rect -1689 762 -1688 772
rect -1662 762 -1661 782
rect -1659 762 -1650 782
rect -1648 762 -1647 782
rect -1624 764 -1623 774
rect -1621 764 -1620 774
rect -2152 709 -2151 729
rect -2149 709 -2141 729
rect -2139 709 -2136 729
rect -2120 714 -2119 724
rect -2117 714 -2101 724
rect -2084 714 -2082 724
rect -2080 714 -2065 724
rect -2035 715 -2034 725
rect -2032 715 -2031 725
rect -1701 691 -1698 701
rect -1695 691 -1692 701
rect -1687 691 -1684 701
rect -1681 691 -1675 701
rect -1646 674 -1645 684
rect -1643 674 -1642 684
rect -1358 621 -1355 631
rect -1352 621 -1349 631
rect -1344 621 -1341 631
rect -1338 621 -1332 631
rect -2165 584 -2164 604
rect -2162 584 -2154 604
rect -2152 584 -2149 604
rect -2133 589 -2132 599
rect -2130 589 -2114 599
rect -2097 589 -2095 599
rect -2093 589 -2078 599
rect -2048 590 -2047 600
rect -2045 590 -2044 600
rect -1303 604 -1302 614
rect -1300 604 -1299 614
rect -1897 565 -1896 575
rect -1894 565 -1893 575
rect -1864 566 -1863 576
rect -1861 566 -1860 576
rect -1835 567 -1832 577
rect -1829 567 -1826 577
rect -1821 567 -1818 577
rect -1815 567 -1809 577
rect -1749 567 -1746 577
rect -1743 567 -1740 577
rect -1735 567 -1732 577
rect -1729 567 -1723 577
rect -1780 550 -1779 560
rect -1777 550 -1776 560
rect -1694 550 -1693 560
rect -1691 550 -1690 560
rect -1664 550 -1663 570
rect -1661 550 -1652 570
rect -1650 550 -1649 570
rect -1626 552 -1625 562
rect -1623 552 -1622 562
rect -1362 520 -1359 530
rect -1356 520 -1353 530
rect -1348 520 -1345 530
rect -1342 520 -1336 530
rect -1331 520 -1330 530
rect -1327 520 -1324 530
rect -1703 479 -1700 489
rect -1697 479 -1694 489
rect -1689 479 -1686 489
rect -1683 479 -1677 489
rect -2165 445 -2164 465
rect -2162 445 -2154 465
rect -2152 445 -2149 465
rect -2133 450 -2132 460
rect -2130 450 -2114 460
rect -2097 450 -2095 460
rect -2093 450 -2078 460
rect -2048 451 -2047 461
rect -2045 451 -2044 461
rect -1230 508 -1229 548
rect -1227 508 -1218 548
rect -1216 508 -1207 548
rect -1205 508 -1197 548
rect -1195 508 -1194 548
rect -1164 518 -1163 528
rect -1161 518 -1160 528
rect -1299 498 -1298 508
rect -1296 498 -1295 508
rect -1648 462 -1647 472
rect -1645 462 -1644 472
rect -540 462 -539 482
rect -537 462 -529 482
rect -527 462 -524 482
rect -508 467 -507 477
rect -505 467 -489 477
rect -472 467 -470 477
rect -468 467 -453 477
rect -423 468 -422 478
rect -420 468 -419 478
rect -1365 398 -1362 408
rect -1359 398 -1356 408
rect -1351 398 -1348 408
rect -1345 398 -1343 408
rect -1339 398 -1337 408
rect -1334 398 -1333 408
rect -1329 398 -1328 408
rect -1325 398 -1323 408
rect -2173 337 -2172 357
rect -2170 337 -2162 357
rect -2160 337 -2157 357
rect -2141 342 -2140 352
rect -2138 342 -2122 352
rect -2105 342 -2103 352
rect -2101 342 -2086 352
rect -2056 343 -2055 353
rect -2053 343 -2052 353
rect -1898 350 -1897 360
rect -1895 350 -1894 360
rect -1865 351 -1864 361
rect -1862 351 -1861 361
rect -1836 352 -1833 362
rect -1830 352 -1827 362
rect -1822 352 -1819 362
rect -1816 352 -1810 362
rect -1750 352 -1747 362
rect -1744 352 -1741 362
rect -1736 352 -1733 362
rect -1730 352 -1724 362
rect -1781 335 -1780 345
rect -1778 335 -1777 345
rect -1695 335 -1694 345
rect -1692 335 -1691 345
rect -1665 335 -1664 355
rect -1662 335 -1653 355
rect -1651 335 -1650 355
rect -1302 376 -1301 386
rect -1299 376 -1298 386
rect -1007 379 -1006 389
rect -1004 379 -1003 389
rect -974 380 -973 390
rect -971 380 -970 390
rect -945 381 -942 391
rect -939 381 -936 391
rect -931 381 -928 391
rect -925 381 -919 391
rect -859 381 -856 391
rect -853 381 -850 391
rect -845 381 -842 391
rect -839 381 -833 391
rect -1627 337 -1626 347
rect -1624 337 -1623 347
rect -890 364 -889 374
rect -887 364 -886 374
rect -804 364 -803 374
rect -801 364 -800 374
rect -774 364 -773 384
rect -771 364 -762 384
rect -760 364 -759 384
rect -736 366 -735 376
rect -733 366 -732 376
rect -538 361 -537 381
rect -535 361 -527 381
rect -525 361 -522 381
rect -506 366 -505 376
rect -503 366 -487 376
rect -470 366 -468 376
rect -466 366 -451 376
rect -421 367 -420 377
rect -418 367 -417 377
rect -1704 264 -1701 274
rect -1698 264 -1695 274
rect -1690 264 -1687 274
rect -1684 264 -1678 274
rect -1376 264 -1373 274
rect -1370 264 -1367 274
rect -1362 264 -1359 274
rect -1356 264 -1350 274
rect -2179 228 -2178 248
rect -2176 228 -2168 248
rect -2166 228 -2163 248
rect -2147 233 -2146 243
rect -2144 233 -2128 243
rect -2111 233 -2109 243
rect -2107 233 -2092 243
rect -2062 234 -2061 244
rect -2059 234 -2058 244
rect -1649 247 -1648 257
rect -1646 247 -1645 257
rect -1007 262 -1006 272
rect -1004 262 -1003 272
rect -974 263 -973 273
rect -971 263 -970 273
rect -945 264 -942 274
rect -939 264 -936 274
rect -931 264 -928 274
rect -925 264 -919 274
rect -859 264 -856 274
rect -853 264 -850 274
rect -845 264 -842 274
rect -839 264 -833 274
rect -1321 247 -1320 257
rect -1318 247 -1317 257
rect -1269 215 -1268 245
rect -1266 215 -1257 245
rect -1255 215 -1244 245
rect -1242 215 -1233 245
rect -1203 224 -1202 234
rect -1200 224 -1199 234
rect -890 247 -889 257
rect -887 247 -886 257
rect -804 247 -803 257
rect -801 247 -800 257
rect -774 247 -773 267
rect -771 247 -762 267
rect -760 247 -759 267
rect -736 249 -735 259
rect -733 249 -732 259
rect -551 236 -550 256
rect -548 236 -540 256
rect -538 236 -535 256
rect -519 241 -518 251
rect -516 241 -500 251
rect -483 241 -481 251
rect -479 241 -464 251
rect -434 242 -433 252
rect -431 242 -430 252
rect -1380 163 -1377 173
rect -1374 163 -1371 173
rect -1366 163 -1363 173
rect -1360 163 -1354 173
rect -1349 163 -1348 173
rect -1345 163 -1342 173
rect -1895 122 -1894 132
rect -1892 122 -1891 132
rect -1862 123 -1861 133
rect -1859 123 -1858 133
rect -1833 124 -1830 134
rect -1827 124 -1824 134
rect -1819 124 -1816 134
rect -1813 124 -1807 134
rect -1747 124 -1744 134
rect -1741 124 -1738 134
rect -1733 124 -1730 134
rect -1727 124 -1721 134
rect -2173 100 -2172 120
rect -2170 100 -2162 120
rect -2160 100 -2157 120
rect -2141 105 -2140 115
rect -2138 105 -2122 115
rect -2105 105 -2103 115
rect -2101 105 -2086 115
rect -2056 106 -2055 116
rect -2053 106 -2052 116
rect -1778 107 -1777 117
rect -1775 107 -1774 117
rect -1692 107 -1691 117
rect -1689 107 -1688 117
rect -1662 107 -1661 127
rect -1659 107 -1650 127
rect -1648 107 -1647 127
rect -1624 109 -1623 119
rect -1621 109 -1620 119
rect -1317 141 -1316 151
rect -1314 141 -1313 151
rect -1009 142 -1008 152
rect -1006 142 -1005 152
rect -976 143 -975 153
rect -973 143 -972 153
rect -947 144 -944 154
rect -941 144 -938 154
rect -933 144 -930 154
rect -927 144 -921 154
rect -861 144 -858 154
rect -855 144 -852 154
rect -847 144 -844 154
rect -841 144 -835 154
rect -892 127 -891 137
rect -889 127 -888 137
rect -806 127 -805 137
rect -803 127 -802 137
rect -776 127 -775 147
rect -773 127 -764 147
rect -762 127 -761 147
rect -738 129 -737 139
rect -735 129 -734 139
rect -551 97 -550 117
rect -548 97 -540 117
rect -538 97 -535 117
rect -519 102 -518 112
rect -516 102 -500 112
rect -483 102 -481 112
rect -479 102 -464 112
rect -434 103 -433 113
rect -431 103 -430 113
rect -1701 36 -1698 46
rect -1695 36 -1692 46
rect -1687 36 -1684 46
rect -1681 36 -1675 46
rect -1379 43 -1376 53
rect -1373 43 -1370 53
rect -1365 43 -1362 53
rect -1359 43 -1353 53
rect -1646 19 -1645 29
rect -1643 19 -1642 29
rect -1324 26 -1323 36
rect -1321 26 -1320 36
rect -1287 31 -1286 51
rect -1284 31 -1275 51
rect -1273 31 -1272 51
rect -1249 33 -1248 43
rect -1246 33 -1245 43
rect -1009 25 -1008 35
rect -1006 25 -1005 35
rect -976 26 -975 36
rect -973 26 -972 36
rect -947 27 -944 37
rect -941 27 -938 37
rect -933 27 -930 37
rect -927 27 -921 37
rect -861 27 -858 37
rect -855 27 -852 37
rect -847 27 -844 37
rect -841 27 -835 37
rect -892 10 -891 20
rect -889 10 -888 20
rect -806 10 -805 20
rect -803 10 -802 20
rect -776 10 -775 30
rect -773 10 -764 30
rect -762 10 -761 30
rect -738 12 -737 22
rect -735 12 -734 22
rect -559 -11 -558 9
rect -556 -11 -548 9
rect -546 -11 -543 9
rect -527 -6 -526 4
rect -524 -6 -508 4
rect -491 -6 -489 4
rect -487 -6 -472 4
rect -442 -5 -441 5
rect -439 -5 -438 5
rect -2177 -46 -2176 -26
rect -2174 -46 -2166 -26
rect -2164 -46 -2161 -26
rect -2145 -41 -2144 -31
rect -2142 -41 -2126 -31
rect -2109 -41 -2107 -31
rect -2105 -41 -2090 -31
rect -2060 -40 -2059 -30
rect -2057 -40 -2056 -30
rect -2150 -174 -2149 -154
rect -2147 -174 -2139 -154
rect -2137 -174 -2134 -154
rect -2118 -169 -2117 -159
rect -2115 -169 -2099 -159
rect -2082 -169 -2080 -159
rect -2078 -169 -2063 -159
rect -2033 -168 -2032 -158
rect -2030 -168 -2029 -158
<< ndcontact >>
rect -2041 792 -2037 797
rect -2033 792 -2029 797
rect -2158 786 -2154 791
rect -2138 786 -2134 791
rect -2126 781 -2122 791
rect -2103 781 -2099 791
rect -2090 781 -2086 791
rect -2067 781 -2063 791
rect -1899 753 -1895 758
rect -1891 753 -1887 758
rect -1866 754 -1862 759
rect -1858 754 -1854 759
rect -1838 732 -1833 742
rect -1807 732 -1802 742
rect -1782 738 -1778 743
rect -1774 738 -1770 743
rect -1752 732 -1747 742
rect -1721 732 -1716 742
rect -1696 738 -1692 743
rect -1688 738 -1684 743
rect -1628 740 -1624 745
rect -1620 740 -1616 745
rect -1666 733 -1662 738
rect -1657 733 -1653 738
rect -1647 733 -1643 738
rect -2039 691 -2035 696
rect -2031 691 -2027 696
rect -2156 685 -2152 690
rect -2136 685 -2132 690
rect -2124 680 -2120 690
rect -2101 680 -2097 690
rect -2088 680 -2084 690
rect -2065 680 -2061 690
rect -1706 644 -1701 654
rect -1675 644 -1670 654
rect -1650 650 -1646 655
rect -1642 650 -1638 655
rect -2052 566 -2048 571
rect -2044 566 -2040 571
rect -2169 560 -2165 565
rect -2149 560 -2145 565
rect -2137 555 -2133 565
rect -2114 555 -2110 565
rect -2101 555 -2097 565
rect -2078 555 -2074 565
rect -1363 574 -1358 584
rect -1332 574 -1327 584
rect -1307 580 -1303 585
rect -1299 580 -1295 585
rect -1901 541 -1897 546
rect -1893 541 -1889 546
rect -1868 542 -1864 547
rect -1860 542 -1856 547
rect -1840 520 -1835 530
rect -1809 520 -1804 530
rect -1784 526 -1780 531
rect -1776 526 -1772 531
rect -1754 520 -1749 530
rect -1723 520 -1718 530
rect -1698 526 -1694 531
rect -1690 526 -1686 531
rect -1630 528 -1626 533
rect -1622 528 -1618 533
rect -1668 521 -1664 526
rect -1659 521 -1655 526
rect -1649 521 -1645 526
rect -1367 460 -1363 475
rect -1324 460 -1320 475
rect -1303 474 -1299 479
rect -1295 474 -1291 479
rect -1168 494 -1164 499
rect -1160 494 -1156 499
rect -1234 468 -1230 473
rect -1224 468 -1220 473
rect -1212 468 -1208 473
rect -1203 468 -1199 473
rect -1194 468 -1188 473
rect -427 444 -423 449
rect -419 444 -415 449
rect -1708 432 -1703 442
rect -1677 432 -1672 442
rect -1652 438 -1648 443
rect -1644 438 -1640 443
rect -544 438 -540 443
rect -524 438 -520 443
rect -512 433 -508 443
rect -489 433 -485 443
rect -476 433 -472 443
rect -453 433 -449 443
rect -2052 427 -2048 432
rect -2044 427 -2040 432
rect -2169 421 -2165 426
rect -2149 421 -2145 426
rect -2137 416 -2133 426
rect -2114 416 -2110 426
rect -2101 416 -2097 426
rect -2078 416 -2074 426
rect -1902 326 -1898 331
rect -1894 326 -1890 331
rect -1869 327 -1865 332
rect -1861 327 -1857 332
rect -2060 319 -2056 324
rect -2052 319 -2048 324
rect -2177 313 -2173 318
rect -2157 313 -2153 318
rect -2145 308 -2141 318
rect -2122 308 -2118 318
rect -2109 308 -2105 318
rect -2086 308 -2082 318
rect -1841 305 -1836 315
rect -1810 305 -1805 315
rect -1785 311 -1781 316
rect -1777 311 -1773 316
rect -1755 305 -1750 315
rect -1724 305 -1719 315
rect -1699 311 -1695 316
rect -1691 311 -1687 316
rect -1370 333 -1366 353
rect -1322 333 -1318 353
rect -1306 352 -1302 357
rect -1298 352 -1294 357
rect -1011 355 -1007 360
rect -1003 355 -999 360
rect -978 356 -974 361
rect -970 356 -966 361
rect -950 334 -945 344
rect -919 334 -914 344
rect -894 340 -890 345
rect -886 340 -882 345
rect -864 334 -859 344
rect -833 334 -828 344
rect -808 340 -804 345
rect -800 340 -796 345
rect -740 342 -736 347
rect -732 342 -728 347
rect -425 343 -421 348
rect -417 343 -413 348
rect -778 335 -774 340
rect -769 335 -765 340
rect -759 335 -755 340
rect -542 337 -538 342
rect -522 337 -518 342
rect -510 332 -506 342
rect -487 332 -483 342
rect -474 332 -470 342
rect -451 332 -447 342
rect -1631 313 -1627 318
rect -1623 313 -1619 318
rect -1669 306 -1665 311
rect -1660 306 -1656 311
rect -1650 306 -1646 311
rect -1709 217 -1704 227
rect -1678 217 -1673 227
rect -1653 223 -1649 228
rect -1645 223 -1641 228
rect -1381 217 -1376 227
rect -1350 217 -1345 227
rect -1325 223 -1321 228
rect -1317 223 -1313 228
rect -2066 210 -2062 215
rect -2058 210 -2054 215
rect -1011 238 -1007 243
rect -1003 238 -999 243
rect -978 239 -974 244
rect -970 239 -966 244
rect -2183 204 -2179 209
rect -2163 204 -2159 209
rect -2151 199 -2147 209
rect -2128 199 -2124 209
rect -2115 199 -2111 209
rect -2092 199 -2088 209
rect -950 217 -945 227
rect -919 217 -914 227
rect -894 223 -890 228
rect -886 223 -882 228
rect -864 217 -859 227
rect -833 217 -828 227
rect -808 223 -804 228
rect -800 223 -796 228
rect -740 225 -736 230
rect -732 225 -728 230
rect -778 218 -774 223
rect -769 218 -765 223
rect -759 218 -755 223
rect -438 218 -434 223
rect -430 218 -426 223
rect -555 212 -551 217
rect -535 212 -531 217
rect -523 207 -519 217
rect -500 207 -496 217
rect -487 207 -483 217
rect -464 207 -460 217
rect -1207 200 -1203 205
rect -1199 200 -1195 205
rect -1273 176 -1269 180
rect -1263 176 -1259 180
rect -1251 176 -1247 180
rect -1233 176 -1227 180
rect -1899 98 -1895 103
rect -1891 98 -1887 103
rect -1866 99 -1862 104
rect -1858 99 -1854 104
rect -2060 82 -2056 87
rect -2052 82 -2048 87
rect -2177 76 -2173 81
rect -2157 76 -2153 81
rect -2145 71 -2141 81
rect -2122 71 -2118 81
rect -2109 71 -2105 81
rect -2086 71 -2082 81
rect -1838 77 -1833 87
rect -1807 77 -1802 87
rect -1782 83 -1778 88
rect -1774 83 -1770 88
rect -1752 77 -1747 87
rect -1721 77 -1716 87
rect -1696 83 -1692 88
rect -1688 83 -1684 88
rect -1385 103 -1381 118
rect -1342 103 -1338 118
rect -1321 117 -1317 122
rect -1313 117 -1309 122
rect -1013 118 -1009 123
rect -1005 118 -1001 123
rect -980 119 -976 124
rect -972 119 -968 124
rect -952 97 -947 107
rect -921 97 -916 107
rect -896 103 -892 108
rect -888 103 -884 108
rect -866 97 -861 107
rect -835 97 -830 107
rect -810 103 -806 108
rect -802 103 -798 108
rect -742 105 -738 110
rect -734 105 -730 110
rect -780 98 -776 103
rect -771 98 -767 103
rect -761 98 -757 103
rect -1628 85 -1624 90
rect -1620 85 -1616 90
rect -1666 78 -1662 83
rect -1657 78 -1653 83
rect -1647 78 -1643 83
rect -438 79 -434 84
rect -430 79 -426 84
rect -555 73 -551 78
rect -535 73 -531 78
rect -523 68 -519 78
rect -500 68 -496 78
rect -487 68 -483 78
rect -464 68 -460 78
rect -1253 9 -1249 14
rect -1245 9 -1241 14
rect -1706 -11 -1701 -1
rect -1675 -11 -1670 -1
rect -1650 -5 -1646 0
rect -1642 -5 -1638 0
rect -1384 -4 -1379 6
rect -1353 -4 -1348 6
rect -1328 2 -1324 7
rect -1320 2 -1316 7
rect -1291 2 -1287 7
rect -1282 2 -1278 7
rect -1272 2 -1268 7
rect -1013 1 -1009 6
rect -1005 1 -1001 6
rect -980 2 -976 7
rect -972 2 -968 7
rect -952 -20 -947 -10
rect -921 -20 -916 -10
rect -896 -14 -892 -9
rect -888 -14 -884 -9
rect -866 -20 -861 -10
rect -835 -20 -830 -10
rect -810 -14 -806 -9
rect -802 -14 -798 -9
rect -742 -12 -738 -7
rect -734 -12 -730 -7
rect -780 -19 -776 -14
rect -771 -19 -767 -14
rect -761 -19 -757 -14
rect -446 -29 -442 -24
rect -438 -29 -434 -24
rect -563 -35 -559 -30
rect -543 -35 -539 -30
rect -531 -40 -527 -30
rect -508 -40 -504 -30
rect -495 -40 -491 -30
rect -472 -40 -468 -30
rect -2064 -64 -2060 -59
rect -2056 -64 -2052 -59
rect -2181 -70 -2177 -65
rect -2161 -70 -2157 -65
rect -2149 -75 -2145 -65
rect -2126 -75 -2122 -65
rect -2113 -75 -2109 -65
rect -2090 -75 -2086 -65
rect -2037 -192 -2033 -187
rect -2029 -192 -2025 -187
rect -2154 -198 -2150 -193
rect -2134 -198 -2130 -193
rect -2122 -203 -2118 -193
rect -2099 -203 -2095 -193
rect -2086 -203 -2082 -193
rect -2063 -203 -2059 -193
<< pdcontact >>
rect -2158 810 -2154 830
rect -2138 810 -2134 830
rect -2126 815 -2122 825
rect -2103 815 -2099 825
rect -2090 815 -2086 825
rect -2067 815 -2063 825
rect -2041 816 -2037 826
rect -2033 816 -2029 826
rect -1899 777 -1895 787
rect -1891 777 -1887 787
rect -1866 778 -1862 788
rect -1858 778 -1854 788
rect -1838 779 -1833 789
rect -1824 779 -1819 789
rect -1807 779 -1802 789
rect -1752 779 -1747 789
rect -1738 779 -1733 789
rect -1721 779 -1716 789
rect -1782 762 -1778 772
rect -1774 762 -1770 772
rect -1696 762 -1692 772
rect -1688 762 -1684 772
rect -1666 762 -1662 782
rect -1647 762 -1643 782
rect -1628 764 -1624 774
rect -1620 764 -1616 774
rect -2156 709 -2152 729
rect -2136 709 -2132 729
rect -2124 714 -2120 724
rect -2101 714 -2097 724
rect -2088 714 -2084 724
rect -2065 714 -2061 724
rect -2039 715 -2035 725
rect -2031 715 -2027 725
rect -1706 691 -1701 701
rect -1692 691 -1687 701
rect -1675 691 -1670 701
rect -1650 674 -1646 684
rect -1642 674 -1638 684
rect -1363 621 -1358 631
rect -1349 621 -1344 631
rect -1332 621 -1327 631
rect -2169 584 -2165 604
rect -2149 584 -2145 604
rect -2137 589 -2133 599
rect -2114 589 -2110 599
rect -2101 589 -2097 599
rect -2078 589 -2074 599
rect -2052 590 -2048 600
rect -2044 590 -2040 600
rect -1307 604 -1303 614
rect -1299 604 -1295 614
rect -1901 565 -1897 575
rect -1893 565 -1889 575
rect -1868 566 -1864 576
rect -1860 566 -1856 576
rect -1840 567 -1835 577
rect -1826 567 -1821 577
rect -1809 567 -1804 577
rect -1754 567 -1749 577
rect -1740 567 -1735 577
rect -1723 567 -1718 577
rect -1784 550 -1780 560
rect -1776 550 -1772 560
rect -1698 550 -1694 560
rect -1690 550 -1686 560
rect -1668 550 -1664 570
rect -1649 550 -1645 570
rect -1630 552 -1626 562
rect -1622 552 -1618 562
rect -1367 520 -1362 530
rect -1353 520 -1348 530
rect -1336 520 -1331 530
rect -1324 520 -1320 530
rect -1708 479 -1703 489
rect -1694 479 -1689 489
rect -1677 479 -1672 489
rect -2169 445 -2165 465
rect -2149 445 -2145 465
rect -2137 450 -2133 460
rect -2114 450 -2110 460
rect -2101 450 -2097 460
rect -2078 450 -2074 460
rect -2052 451 -2048 461
rect -2044 451 -2040 461
rect -1234 508 -1230 548
rect -1194 508 -1188 548
rect -1168 518 -1164 528
rect -1160 518 -1156 528
rect -1303 498 -1299 508
rect -1295 498 -1291 508
rect -1652 462 -1648 472
rect -1644 462 -1640 472
rect -544 462 -540 482
rect -524 462 -520 482
rect -512 467 -508 477
rect -489 467 -485 477
rect -476 467 -472 477
rect -453 467 -449 477
rect -427 468 -423 478
rect -419 468 -415 478
rect -1370 398 -1365 408
rect -1356 398 -1351 408
rect -1343 398 -1339 408
rect -1333 398 -1329 408
rect -1323 398 -1319 408
rect -2177 337 -2173 357
rect -2157 337 -2153 357
rect -2145 342 -2141 352
rect -2122 342 -2118 352
rect -2109 342 -2105 352
rect -2086 342 -2082 352
rect -2060 343 -2056 353
rect -2052 343 -2048 353
rect -1902 350 -1898 360
rect -1894 350 -1890 360
rect -1869 351 -1865 361
rect -1861 351 -1857 361
rect -1841 352 -1836 362
rect -1827 352 -1822 362
rect -1810 352 -1805 362
rect -1755 352 -1750 362
rect -1741 352 -1736 362
rect -1724 352 -1719 362
rect -1785 335 -1781 345
rect -1777 335 -1773 345
rect -1699 335 -1695 345
rect -1691 335 -1687 345
rect -1669 335 -1665 355
rect -1650 335 -1646 355
rect -1306 376 -1302 386
rect -1298 376 -1294 386
rect -1011 379 -1007 389
rect -1003 379 -999 389
rect -978 380 -974 390
rect -970 380 -966 390
rect -950 381 -945 391
rect -936 381 -931 391
rect -919 381 -914 391
rect -864 381 -859 391
rect -850 381 -845 391
rect -833 381 -828 391
rect -1631 337 -1627 347
rect -1623 337 -1619 347
rect -894 364 -890 374
rect -886 364 -882 374
rect -808 364 -804 374
rect -800 364 -796 374
rect -778 364 -774 384
rect -759 364 -755 384
rect -740 366 -736 376
rect -732 366 -728 376
rect -542 361 -538 381
rect -522 361 -518 381
rect -510 366 -506 376
rect -487 366 -483 376
rect -474 366 -470 376
rect -451 366 -447 376
rect -425 367 -421 377
rect -417 367 -413 377
rect -1709 264 -1704 274
rect -1695 264 -1690 274
rect -1678 264 -1673 274
rect -1381 264 -1376 274
rect -1367 264 -1362 274
rect -1350 264 -1345 274
rect -2183 228 -2179 248
rect -2163 228 -2159 248
rect -2151 233 -2147 243
rect -2128 233 -2124 243
rect -2115 233 -2111 243
rect -2092 233 -2088 243
rect -2066 234 -2062 244
rect -2058 234 -2054 244
rect -1653 247 -1649 257
rect -1645 247 -1641 257
rect -1011 262 -1007 272
rect -1003 262 -999 272
rect -978 263 -974 273
rect -970 263 -966 273
rect -950 264 -945 274
rect -936 264 -931 274
rect -919 264 -914 274
rect -864 264 -859 274
rect -850 264 -845 274
rect -833 264 -828 274
rect -1325 247 -1321 257
rect -1317 247 -1313 257
rect -1273 215 -1269 245
rect -1233 215 -1227 245
rect -1207 224 -1203 234
rect -1199 224 -1195 234
rect -894 247 -890 257
rect -886 247 -882 257
rect -808 247 -804 257
rect -800 247 -796 257
rect -778 247 -774 267
rect -759 247 -755 267
rect -740 249 -736 259
rect -732 249 -728 259
rect -555 236 -551 256
rect -535 236 -531 256
rect -523 241 -519 251
rect -500 241 -496 251
rect -487 241 -483 251
rect -464 241 -460 251
rect -438 242 -434 252
rect -430 242 -426 252
rect -1385 163 -1380 173
rect -1371 163 -1366 173
rect -1354 163 -1349 173
rect -1342 163 -1338 173
rect -1899 122 -1895 132
rect -1891 122 -1887 132
rect -1866 123 -1862 133
rect -1858 123 -1854 133
rect -1838 124 -1833 134
rect -1824 124 -1819 134
rect -1807 124 -1802 134
rect -1752 124 -1747 134
rect -1738 124 -1733 134
rect -1721 124 -1716 134
rect -2177 100 -2173 120
rect -2157 100 -2153 120
rect -2145 105 -2141 115
rect -2122 105 -2118 115
rect -2109 105 -2105 115
rect -2086 105 -2082 115
rect -2060 106 -2056 116
rect -2052 106 -2048 116
rect -1782 107 -1778 117
rect -1774 107 -1770 117
rect -1696 107 -1692 117
rect -1688 107 -1684 117
rect -1666 107 -1662 127
rect -1647 107 -1643 127
rect -1628 109 -1624 119
rect -1620 109 -1616 119
rect -1321 141 -1317 151
rect -1313 141 -1309 151
rect -1013 142 -1009 152
rect -1005 142 -1001 152
rect -980 143 -976 153
rect -972 143 -968 153
rect -952 144 -947 154
rect -938 144 -933 154
rect -921 144 -916 154
rect -866 144 -861 154
rect -852 144 -847 154
rect -835 144 -830 154
rect -896 127 -892 137
rect -888 127 -884 137
rect -810 127 -806 137
rect -802 127 -798 137
rect -780 127 -776 147
rect -761 127 -757 147
rect -742 129 -738 139
rect -734 129 -730 139
rect -555 97 -551 117
rect -535 97 -531 117
rect -523 102 -519 112
rect -500 102 -496 112
rect -487 102 -483 112
rect -464 102 -460 112
rect -438 103 -434 113
rect -430 103 -426 113
rect -1706 36 -1701 46
rect -1692 36 -1687 46
rect -1675 36 -1670 46
rect -1384 43 -1379 53
rect -1370 43 -1365 53
rect -1353 43 -1348 53
rect -1650 19 -1646 29
rect -1642 19 -1638 29
rect -1328 26 -1324 36
rect -1320 26 -1316 36
rect -1291 31 -1287 51
rect -1272 31 -1268 51
rect -1253 33 -1249 43
rect -1245 33 -1241 43
rect -1013 25 -1009 35
rect -1005 25 -1001 35
rect -980 26 -976 36
rect -972 26 -968 36
rect -952 27 -947 37
rect -938 27 -933 37
rect -921 27 -916 37
rect -866 27 -861 37
rect -852 27 -847 37
rect -835 27 -830 37
rect -896 10 -892 20
rect -888 10 -884 20
rect -810 10 -806 20
rect -802 10 -798 20
rect -780 10 -776 30
rect -761 10 -757 30
rect -742 12 -738 22
rect -734 12 -730 22
rect -563 -11 -559 9
rect -543 -11 -539 9
rect -531 -6 -527 4
rect -508 -6 -504 4
rect -495 -6 -491 4
rect -472 -6 -468 4
rect -446 -5 -442 5
rect -438 -5 -434 5
rect -2181 -46 -2177 -26
rect -2161 -46 -2157 -26
rect -2149 -41 -2145 -31
rect -2126 -41 -2122 -31
rect -2113 -41 -2109 -31
rect -2090 -41 -2086 -31
rect -2064 -40 -2060 -30
rect -2056 -40 -2052 -30
rect -2154 -174 -2150 -154
rect -2134 -174 -2130 -154
rect -2122 -169 -2118 -159
rect -2099 -169 -2095 -159
rect -2086 -169 -2082 -159
rect -2063 -169 -2059 -159
rect -2037 -168 -2033 -158
rect -2029 -168 -2025 -158
<< polysilicon >>
rect -2153 830 -2151 833
rect -2143 830 -2141 833
rect -2121 825 -2119 829
rect -2084 825 -2082 829
rect -2036 826 -2034 830
rect -2153 791 -2151 810
rect -2143 794 -2141 810
rect -2121 791 -2119 815
rect -2110 791 -2108 798
rect -2084 791 -2082 815
rect -2073 791 -2071 798
rect -2036 797 -2034 816
rect -2153 783 -2151 786
rect -2036 786 -2034 792
rect -1894 787 -1892 791
rect -1861 788 -1859 792
rect -1830 789 -1827 793
rect -1816 789 -1813 793
rect -1744 789 -1741 793
rect -1730 789 -1727 793
rect -2121 778 -2119 781
rect -2110 778 -2108 781
rect -2084 778 -2082 781
rect -2073 778 -2071 781
rect -1661 782 -1659 785
rect -1650 782 -1648 785
rect -1894 758 -1892 777
rect -1861 759 -1859 778
rect -1830 759 -1827 779
rect -1894 747 -1892 753
rect -1861 748 -1859 754
rect -1830 742 -1827 754
rect -1816 751 -1813 779
rect -1777 772 -1775 776
rect -1816 742 -1813 746
rect -1777 743 -1775 762
rect -1744 759 -1741 779
rect -1744 742 -1741 754
rect -1730 751 -1727 779
rect -1691 772 -1689 776
rect -1623 774 -1621 778
rect -1730 742 -1727 746
rect -1691 743 -1689 762
rect -1777 732 -1775 738
rect -1661 738 -1659 762
rect -1650 738 -1648 762
rect -1623 745 -1621 764
rect -1691 732 -1689 738
rect -1623 734 -1621 740
rect -2151 729 -2149 732
rect -2141 729 -2139 732
rect -1830 729 -1827 732
rect -1816 729 -1813 732
rect -1744 729 -1741 732
rect -1730 729 -1727 732
rect -1661 730 -1659 733
rect -1650 730 -1648 733
rect -2119 724 -2117 728
rect -2082 724 -2080 728
rect -2034 725 -2032 729
rect -2151 690 -2149 709
rect -2141 693 -2139 709
rect -2119 690 -2117 714
rect -2108 690 -2106 697
rect -2082 690 -2080 714
rect -2071 690 -2069 697
rect -2034 696 -2032 715
rect -1698 701 -1695 705
rect -1684 701 -1681 705
rect -2151 682 -2149 685
rect -2034 685 -2032 691
rect -2119 677 -2117 680
rect -2108 677 -2106 680
rect -2082 677 -2080 680
rect -2071 677 -2069 680
rect -1698 671 -1695 691
rect -1698 654 -1695 666
rect -1684 663 -1681 691
rect -1645 684 -1643 688
rect -1684 654 -1681 658
rect -1645 655 -1643 674
rect -1645 644 -1643 650
rect -1698 641 -1695 644
rect -1684 641 -1681 644
rect -1355 631 -1352 635
rect -1341 631 -1338 635
rect -2164 604 -2162 607
rect -2154 604 -2152 607
rect -2132 599 -2130 603
rect -2095 599 -2093 603
rect -2047 600 -2045 604
rect -1355 601 -1352 621
rect -2164 565 -2162 584
rect -2154 568 -2152 584
rect -2132 565 -2130 589
rect -2121 565 -2119 572
rect -2095 565 -2093 589
rect -2084 565 -2082 572
rect -2047 571 -2045 590
rect -1355 584 -1352 596
rect -1341 593 -1338 621
rect -1302 614 -1300 618
rect -1341 584 -1338 588
rect -1302 585 -1300 604
rect -1896 575 -1894 579
rect -1863 576 -1861 580
rect -1832 577 -1829 581
rect -1818 577 -1815 581
rect -1746 577 -1743 581
rect -1732 577 -1729 581
rect -2164 557 -2162 560
rect -2047 560 -2045 566
rect -1302 574 -1300 580
rect -1663 570 -1661 573
rect -1652 570 -1650 573
rect -1355 571 -1352 574
rect -1341 571 -1338 574
rect -2132 552 -2130 555
rect -2121 552 -2119 555
rect -2095 552 -2093 555
rect -2084 552 -2082 555
rect -1896 546 -1894 565
rect -1863 547 -1861 566
rect -1832 547 -1829 567
rect -1896 535 -1894 541
rect -1863 536 -1861 542
rect -1832 530 -1829 542
rect -1818 539 -1815 567
rect -1779 560 -1777 564
rect -1818 530 -1815 534
rect -1779 531 -1777 550
rect -1746 547 -1743 567
rect -1746 530 -1743 542
rect -1732 539 -1729 567
rect -1693 560 -1691 564
rect -1625 562 -1623 566
rect -1732 530 -1729 534
rect -1693 531 -1691 550
rect -1779 520 -1777 526
rect -1663 526 -1661 550
rect -1652 526 -1650 550
rect -1625 533 -1623 552
rect -1229 548 -1227 551
rect -1218 548 -1216 551
rect -1207 548 -1205 551
rect -1197 548 -1195 551
rect -1359 530 -1356 534
rect -1345 530 -1342 534
rect -1330 530 -1327 534
rect -1693 520 -1691 526
rect -1625 522 -1623 528
rect -1832 517 -1829 520
rect -1818 517 -1815 520
rect -1746 517 -1743 520
rect -1732 517 -1729 520
rect -1663 518 -1661 521
rect -1652 518 -1650 521
rect -1700 489 -1697 493
rect -1686 489 -1683 493
rect -2164 465 -2162 468
rect -2154 465 -2152 468
rect -2132 460 -2130 464
rect -2095 460 -2093 464
rect -2047 461 -2045 465
rect -1700 459 -1697 479
rect -2164 426 -2162 445
rect -2154 429 -2152 445
rect -2132 426 -2130 450
rect -2121 426 -2119 433
rect -2095 426 -2093 450
rect -2084 426 -2082 433
rect -2047 432 -2045 451
rect -1700 442 -1697 454
rect -1686 451 -1683 479
rect -1647 472 -1645 476
rect -1359 475 -1356 520
rect -1345 475 -1342 520
rect -1330 475 -1327 520
rect -1298 508 -1296 512
rect -1163 528 -1161 532
rect -1298 479 -1296 498
rect -1686 442 -1683 446
rect -1647 443 -1645 462
rect -1298 468 -1296 474
rect -1229 473 -1227 508
rect -1218 473 -1216 508
rect -1207 473 -1205 508
rect -1197 473 -1195 508
rect -1163 499 -1161 518
rect -1163 488 -1161 494
rect -539 482 -537 485
rect -529 482 -527 485
rect -1229 465 -1227 468
rect -1218 465 -1216 468
rect -1207 465 -1205 468
rect -1197 465 -1195 468
rect -507 477 -505 481
rect -470 477 -468 481
rect -422 478 -420 482
rect -1359 456 -1356 460
rect -1345 456 -1342 460
rect -1330 456 -1327 460
rect -539 443 -537 462
rect -529 446 -527 462
rect -507 443 -505 467
rect -496 443 -494 450
rect -470 443 -468 467
rect -459 443 -457 450
rect -422 449 -420 468
rect -1647 432 -1645 438
rect -539 435 -537 438
rect -422 438 -420 444
rect -1700 429 -1697 432
rect -1686 429 -1683 432
rect -507 430 -505 433
rect -496 430 -494 433
rect -470 430 -468 433
rect -459 430 -457 433
rect -2164 418 -2162 421
rect -2047 421 -2045 427
rect -2132 413 -2130 416
rect -2121 413 -2119 416
rect -2095 413 -2093 416
rect -2084 413 -2082 416
rect -1362 408 -1359 412
rect -1348 408 -1345 412
rect -1337 408 -1334 412
rect -1328 408 -1325 412
rect -1897 360 -1895 364
rect -1864 361 -1862 365
rect -1833 362 -1830 366
rect -1819 362 -1816 366
rect -1747 362 -1744 366
rect -1733 362 -1730 366
rect -2172 357 -2170 360
rect -2162 357 -2160 360
rect -2140 352 -2138 356
rect -2103 352 -2101 356
rect -2055 353 -2053 357
rect -1664 355 -1662 358
rect -1653 355 -1651 358
rect -2172 318 -2170 337
rect -2162 321 -2160 337
rect -2140 318 -2138 342
rect -2129 318 -2127 325
rect -2103 318 -2101 342
rect -2092 318 -2090 325
rect -2055 324 -2053 343
rect -1897 331 -1895 350
rect -1864 332 -1862 351
rect -1833 332 -1830 352
rect -1897 320 -1895 326
rect -1864 321 -1862 327
rect -2172 310 -2170 313
rect -2055 313 -2053 319
rect -1833 315 -1830 327
rect -1819 324 -1816 352
rect -1780 345 -1778 349
rect -1819 315 -1816 319
rect -1780 316 -1778 335
rect -1747 332 -1744 352
rect -2140 305 -2138 308
rect -2129 305 -2127 308
rect -2103 305 -2101 308
rect -2092 305 -2090 308
rect -1747 315 -1744 327
rect -1733 324 -1730 352
rect -1694 345 -1692 349
rect -1362 353 -1359 398
rect -1348 353 -1345 398
rect -1337 364 -1334 398
rect -1336 359 -1334 364
rect -1328 359 -1325 398
rect -1301 386 -1299 390
rect -1006 389 -1004 393
rect -973 390 -971 394
rect -942 391 -939 395
rect -928 391 -925 395
rect -856 391 -853 395
rect -842 391 -839 395
rect -773 384 -771 387
rect -762 384 -760 387
rect -1337 353 -1334 359
rect -1301 357 -1299 376
rect -1006 360 -1004 379
rect -973 361 -971 380
rect -942 361 -939 381
rect -1328 353 -1325 354
rect -1626 347 -1624 351
rect -1733 315 -1730 319
rect -1694 316 -1692 335
rect -1780 305 -1778 311
rect -1664 311 -1662 335
rect -1653 311 -1651 335
rect -1626 318 -1624 337
rect -1301 346 -1299 352
rect -1006 349 -1004 355
rect -973 350 -971 356
rect -942 344 -939 356
rect -928 353 -925 381
rect -889 374 -887 378
rect -928 344 -925 348
rect -889 345 -887 364
rect -856 361 -853 381
rect -856 344 -853 356
rect -842 353 -839 381
rect -803 374 -801 378
rect -537 381 -535 384
rect -527 381 -525 384
rect -735 376 -733 380
rect -842 344 -839 348
rect -803 345 -801 364
rect -889 334 -887 340
rect -773 340 -771 364
rect -762 340 -760 364
rect -735 347 -733 366
rect -505 376 -503 380
rect -468 376 -466 380
rect -420 377 -418 381
rect -537 342 -535 361
rect -527 345 -525 361
rect -505 342 -503 366
rect -494 342 -492 349
rect -468 342 -466 366
rect -457 342 -455 349
rect -420 348 -418 367
rect -803 334 -801 340
rect -735 336 -733 342
rect -1362 330 -1359 333
rect -1348 330 -1345 333
rect -1337 330 -1334 333
rect -1328 330 -1325 333
rect -942 331 -939 334
rect -928 331 -925 334
rect -856 331 -853 334
rect -842 331 -839 334
rect -773 332 -771 335
rect -762 332 -760 335
rect -537 334 -535 337
rect -420 337 -418 343
rect -505 329 -503 332
rect -494 329 -492 332
rect -468 329 -466 332
rect -457 329 -455 332
rect -1694 305 -1692 311
rect -1626 307 -1624 313
rect -1833 302 -1830 305
rect -1819 302 -1816 305
rect -1747 302 -1744 305
rect -1733 302 -1730 305
rect -1664 303 -1662 306
rect -1653 303 -1651 306
rect -1701 274 -1698 278
rect -1687 274 -1684 278
rect -1373 274 -1370 278
rect -1359 274 -1356 278
rect -1006 272 -1004 276
rect -973 273 -971 277
rect -942 274 -939 278
rect -928 274 -925 278
rect -856 274 -853 278
rect -842 274 -839 278
rect -2178 248 -2176 251
rect -2168 248 -2166 251
rect -2146 243 -2144 247
rect -2109 243 -2107 247
rect -2061 244 -2059 248
rect -1701 244 -1698 264
rect -2178 209 -2176 228
rect -2168 212 -2166 228
rect -2146 209 -2144 233
rect -2135 209 -2133 216
rect -2109 209 -2107 233
rect -2098 209 -2096 216
rect -2061 215 -2059 234
rect -1701 227 -1698 239
rect -1687 236 -1684 264
rect -1648 257 -1646 261
rect -1687 227 -1684 231
rect -1648 228 -1646 247
rect -1373 244 -1370 264
rect -1373 227 -1370 239
rect -1359 236 -1356 264
rect -773 267 -771 270
rect -762 267 -760 270
rect -1320 257 -1318 261
rect -1359 227 -1356 231
rect -1320 228 -1318 247
rect -1268 245 -1266 250
rect -1257 245 -1255 250
rect -1244 245 -1242 250
rect -1648 217 -1646 223
rect -1320 217 -1318 223
rect -1701 214 -1698 217
rect -1687 214 -1684 217
rect -1373 214 -1370 217
rect -1359 214 -1356 217
rect -1006 243 -1004 262
rect -973 244 -971 263
rect -942 244 -939 264
rect -1202 234 -1200 238
rect -1006 232 -1004 238
rect -973 233 -971 239
rect -942 227 -939 239
rect -928 236 -925 264
rect -889 257 -887 261
rect -928 227 -925 231
rect -889 228 -887 247
rect -856 244 -853 264
rect -2178 201 -2176 204
rect -2061 204 -2059 210
rect -2146 196 -2144 199
rect -2135 196 -2133 199
rect -2109 196 -2107 199
rect -2098 196 -2096 199
rect -1268 180 -1266 215
rect -1257 180 -1255 215
rect -1244 180 -1242 215
rect -1202 205 -1200 224
rect -856 227 -853 239
rect -842 236 -839 264
rect -803 257 -801 261
rect -735 259 -733 263
rect -550 256 -548 259
rect -540 256 -538 259
rect -842 227 -839 231
rect -803 228 -801 247
rect -889 217 -887 223
rect -773 223 -771 247
rect -762 223 -760 247
rect -735 230 -733 249
rect -518 251 -516 255
rect -481 251 -479 255
rect -433 252 -431 256
rect -803 217 -801 223
rect -735 219 -733 225
rect -942 214 -939 217
rect -928 214 -925 217
rect -856 214 -853 217
rect -842 214 -839 217
rect -773 215 -771 218
rect -762 215 -760 218
rect -550 217 -548 236
rect -540 220 -538 236
rect -518 217 -516 241
rect -507 217 -505 224
rect -481 217 -479 241
rect -470 217 -468 224
rect -433 223 -431 242
rect -550 209 -548 212
rect -433 212 -431 218
rect -518 204 -516 207
rect -507 204 -505 207
rect -481 204 -479 207
rect -470 204 -468 207
rect -1202 194 -1200 200
rect -1377 173 -1374 177
rect -1363 173 -1360 177
rect -1348 173 -1345 177
rect -1268 173 -1266 176
rect -1257 173 -1255 176
rect -1244 173 -1242 176
rect -1894 132 -1892 136
rect -1861 133 -1859 137
rect -1830 134 -1827 138
rect -1816 134 -1813 138
rect -1744 134 -1741 138
rect -1730 134 -1727 138
rect -2172 120 -2170 123
rect -2162 120 -2160 123
rect -1661 127 -1659 130
rect -1650 127 -1648 130
rect -2140 115 -2138 119
rect -2103 115 -2101 119
rect -2055 116 -2053 120
rect -2172 81 -2170 100
rect -2162 84 -2160 100
rect -2140 81 -2138 105
rect -2129 81 -2127 88
rect -2103 81 -2101 105
rect -2092 81 -2090 88
rect -2055 87 -2053 106
rect -1894 103 -1892 122
rect -1861 104 -1859 123
rect -1830 104 -1827 124
rect -1894 92 -1892 98
rect -1861 93 -1859 99
rect -1830 87 -1827 99
rect -1816 96 -1813 124
rect -1777 117 -1775 121
rect -1816 87 -1813 91
rect -1777 88 -1775 107
rect -1744 104 -1741 124
rect -2172 73 -2170 76
rect -2055 76 -2053 82
rect -1744 87 -1741 99
rect -1730 96 -1727 124
rect -1691 117 -1689 121
rect -1623 119 -1621 123
rect -1377 118 -1374 163
rect -1363 118 -1360 163
rect -1348 118 -1345 163
rect -1316 151 -1314 155
rect -1008 152 -1006 156
rect -975 153 -973 157
rect -944 154 -941 158
rect -930 154 -927 158
rect -858 154 -855 158
rect -844 154 -841 158
rect -775 147 -773 150
rect -764 147 -762 150
rect -1316 122 -1314 141
rect -1008 123 -1006 142
rect -975 124 -973 143
rect -944 124 -941 144
rect -1730 87 -1727 91
rect -1691 88 -1689 107
rect -1777 77 -1775 83
rect -1661 83 -1659 107
rect -1650 83 -1648 107
rect -1623 90 -1621 109
rect -1316 111 -1314 117
rect -1008 112 -1006 118
rect -975 113 -973 119
rect -944 107 -941 119
rect -930 116 -927 144
rect -891 137 -889 141
rect -930 107 -927 111
rect -891 108 -889 127
rect -858 124 -855 144
rect -1377 99 -1374 103
rect -1363 99 -1360 103
rect -1348 99 -1345 103
rect -858 107 -855 119
rect -844 116 -841 144
rect -805 137 -803 141
rect -737 139 -735 143
rect -844 107 -841 111
rect -805 108 -803 127
rect -891 97 -889 103
rect -775 103 -773 127
rect -764 103 -762 127
rect -737 110 -735 129
rect -550 117 -548 120
rect -540 117 -538 120
rect -805 97 -803 103
rect -737 99 -735 105
rect -944 94 -941 97
rect -930 94 -927 97
rect -858 94 -855 97
rect -844 94 -841 97
rect -775 95 -773 98
rect -764 95 -762 98
rect -518 112 -516 116
rect -481 112 -479 116
rect -433 113 -431 117
rect -1691 77 -1689 83
rect -1623 79 -1621 85
rect -550 78 -548 97
rect -540 81 -538 97
rect -518 78 -516 102
rect -507 78 -505 85
rect -481 78 -479 102
rect -470 78 -468 85
rect -433 84 -431 103
rect -1830 74 -1827 77
rect -1816 74 -1813 77
rect -1744 74 -1741 77
rect -1730 74 -1727 77
rect -1661 75 -1659 78
rect -1650 75 -1648 78
rect -2140 68 -2138 71
rect -2129 68 -2127 71
rect -2103 68 -2101 71
rect -2092 68 -2090 71
rect -550 70 -548 73
rect -433 73 -431 79
rect -518 65 -516 68
rect -507 65 -505 68
rect -481 65 -479 68
rect -470 65 -468 68
rect -1376 53 -1373 57
rect -1362 53 -1359 57
rect -1698 46 -1695 50
rect -1684 46 -1681 50
rect -1286 51 -1284 54
rect -1275 51 -1273 54
rect -1698 16 -1695 36
rect -1698 -1 -1695 11
rect -1684 8 -1681 36
rect -1645 29 -1643 33
rect -1376 23 -1373 43
rect -1684 -1 -1681 3
rect -1645 0 -1643 19
rect -1376 6 -1373 18
rect -1362 15 -1359 43
rect -1323 36 -1321 40
rect -1248 43 -1246 47
rect -1008 35 -1006 39
rect -975 36 -973 40
rect -944 37 -941 41
rect -930 37 -927 41
rect -858 37 -855 41
rect -844 37 -841 41
rect -1362 6 -1359 10
rect -1323 7 -1321 26
rect -1286 7 -1284 31
rect -1275 7 -1273 31
rect -1248 14 -1246 33
rect -775 30 -773 33
rect -764 30 -762 33
rect -1248 3 -1246 9
rect -1008 6 -1006 25
rect -975 7 -973 26
rect -944 7 -941 27
rect -1323 -4 -1321 2
rect -1286 -1 -1284 2
rect -1275 -1 -1273 2
rect -1645 -11 -1643 -5
rect -1376 -7 -1373 -4
rect -1362 -7 -1359 -4
rect -1008 -5 -1006 1
rect -975 -4 -973 2
rect -944 -10 -941 2
rect -930 -1 -927 27
rect -891 20 -889 24
rect -930 -10 -927 -6
rect -891 -9 -889 10
rect -858 7 -855 27
rect -1698 -14 -1695 -11
rect -1684 -14 -1681 -11
rect -858 -10 -855 2
rect -844 -1 -841 27
rect -805 20 -803 24
rect -737 22 -735 26
rect -844 -10 -841 -6
rect -805 -9 -803 10
rect -891 -20 -889 -14
rect -775 -14 -773 10
rect -764 -14 -762 10
rect -737 -7 -735 12
rect -558 9 -556 12
rect -548 9 -546 12
rect -526 4 -524 8
rect -489 4 -487 8
rect -441 5 -439 9
rect -805 -20 -803 -14
rect -737 -18 -735 -12
rect -944 -23 -941 -20
rect -930 -23 -927 -20
rect -858 -23 -855 -20
rect -844 -23 -841 -20
rect -775 -22 -773 -19
rect -764 -22 -762 -19
rect -2176 -26 -2174 -23
rect -2166 -26 -2164 -23
rect -2144 -31 -2142 -27
rect -2107 -31 -2105 -27
rect -2059 -30 -2057 -26
rect -558 -30 -556 -11
rect -548 -27 -546 -11
rect -526 -30 -524 -6
rect -515 -30 -513 -23
rect -489 -30 -487 -6
rect -478 -30 -476 -23
rect -441 -24 -439 -5
rect -558 -38 -556 -35
rect -441 -35 -439 -29
rect -2176 -65 -2174 -46
rect -2166 -62 -2164 -46
rect -2144 -65 -2142 -41
rect -2133 -65 -2131 -58
rect -2107 -65 -2105 -41
rect -2096 -65 -2094 -58
rect -2059 -59 -2057 -40
rect -526 -43 -524 -40
rect -515 -43 -513 -40
rect -489 -43 -487 -40
rect -478 -43 -476 -40
rect -2176 -73 -2174 -70
rect -2059 -70 -2057 -64
rect -2144 -78 -2142 -75
rect -2133 -78 -2131 -75
rect -2107 -78 -2105 -75
rect -2096 -78 -2094 -75
rect -2149 -154 -2147 -151
rect -2139 -154 -2137 -151
rect -2117 -159 -2115 -155
rect -2080 -159 -2078 -155
rect -2032 -158 -2030 -154
rect -2149 -193 -2147 -174
rect -2139 -190 -2137 -174
rect -2117 -193 -2115 -169
rect -2106 -193 -2104 -186
rect -2080 -193 -2078 -169
rect -2069 -193 -2067 -186
rect -2032 -187 -2030 -168
rect -2149 -201 -2147 -198
rect -2032 -198 -2030 -192
rect -2117 -206 -2115 -203
rect -2106 -206 -2104 -203
rect -2080 -206 -2078 -203
rect -2069 -206 -2067 -203
<< polycontact >>
rect -2157 798 -2153 802
rect -2147 794 -2143 798
rect -2125 798 -2121 802
rect -2088 798 -2084 802
rect -2114 794 -2110 798
rect -2040 800 -2036 804
rect -2077 794 -2073 798
rect -1898 761 -1894 765
rect -1865 762 -1861 766
rect -1832 754 -1827 759
rect -1818 746 -1813 751
rect -1781 746 -1777 750
rect -1746 754 -1741 759
rect -1732 746 -1727 751
rect -1695 746 -1691 750
rect -1665 749 -1661 753
rect -1654 749 -1650 753
rect -1627 748 -1623 752
rect -2155 697 -2151 701
rect -2145 693 -2141 697
rect -2123 697 -2119 701
rect -2086 697 -2082 701
rect -2112 693 -2108 697
rect -2038 699 -2034 703
rect -2075 693 -2071 697
rect -1700 666 -1695 671
rect -1686 658 -1681 663
rect -1649 658 -1645 662
rect -1357 596 -1352 601
rect -2168 572 -2164 576
rect -2158 568 -2154 572
rect -2136 572 -2132 576
rect -2099 572 -2095 576
rect -2125 568 -2121 572
rect -2051 574 -2047 578
rect -2088 568 -2084 572
rect -1343 588 -1338 593
rect -1306 588 -1302 592
rect -1900 549 -1896 553
rect -1867 550 -1863 554
rect -1834 542 -1829 547
rect -1820 534 -1815 539
rect -1783 534 -1779 538
rect -1748 542 -1743 547
rect -1734 534 -1729 539
rect -1697 534 -1693 538
rect -1667 537 -1663 541
rect -1656 537 -1652 541
rect -1629 536 -1625 540
rect -1364 495 -1359 500
rect -1702 454 -1697 459
rect -2168 433 -2164 437
rect -2158 429 -2154 433
rect -2136 433 -2132 437
rect -2099 433 -2095 437
rect -2125 429 -2121 433
rect -2051 435 -2047 439
rect -2088 429 -2084 433
rect -1350 487 -1345 492
rect -1335 478 -1330 483
rect -1302 482 -1298 486
rect -1233 496 -1229 500
rect -1688 446 -1683 451
rect -1651 446 -1647 450
rect -1222 489 -1218 493
rect -1211 482 -1207 486
rect -1201 483 -1197 487
rect -1167 502 -1163 506
rect -543 450 -539 454
rect -533 446 -529 450
rect -511 450 -507 454
rect -474 450 -470 454
rect -500 446 -496 450
rect -426 452 -422 456
rect -463 446 -459 450
rect -1367 373 -1362 378
rect -2176 325 -2172 329
rect -2166 321 -2162 325
rect -2144 325 -2140 329
rect -2107 325 -2103 329
rect -2133 321 -2129 325
rect -2059 327 -2055 331
rect -2096 321 -2092 325
rect -1901 334 -1897 338
rect -1868 335 -1864 339
rect -1835 327 -1830 332
rect -1821 319 -1816 324
rect -1784 319 -1780 323
rect -1749 327 -1744 332
rect -1353 365 -1348 370
rect -1341 359 -1336 364
rect -1305 360 -1301 364
rect -1330 354 -1325 359
rect -1010 363 -1006 367
rect -977 364 -973 368
rect -1735 319 -1730 324
rect -1698 319 -1694 323
rect -1668 322 -1664 326
rect -1657 322 -1653 326
rect -1630 321 -1626 325
rect -944 356 -939 361
rect -930 348 -925 353
rect -893 348 -889 352
rect -858 356 -853 361
rect -844 348 -839 353
rect -807 348 -803 352
rect -777 351 -773 355
rect -766 351 -762 355
rect -739 350 -735 354
rect -541 349 -537 353
rect -531 345 -527 349
rect -509 349 -505 353
rect -472 349 -468 353
rect -498 345 -494 349
rect -424 351 -420 355
rect -461 345 -457 349
rect -1703 239 -1698 244
rect -2182 216 -2178 220
rect -2172 212 -2168 216
rect -2150 216 -2146 220
rect -2113 216 -2109 220
rect -2139 212 -2135 216
rect -2065 218 -2061 222
rect -2102 212 -2098 216
rect -1689 231 -1684 236
rect -1652 231 -1648 235
rect -1375 239 -1370 244
rect -1361 231 -1356 236
rect -1324 231 -1320 235
rect -1010 246 -1006 250
rect -977 247 -973 251
rect -944 239 -939 244
rect -930 231 -925 236
rect -893 231 -889 235
rect -858 239 -853 244
rect -1272 202 -1268 206
rect -1261 196 -1257 200
rect -1248 189 -1244 193
rect -1206 208 -1202 212
rect -844 231 -839 236
rect -807 231 -803 235
rect -777 234 -773 238
rect -766 234 -762 238
rect -739 233 -735 237
rect -554 224 -550 228
rect -544 220 -540 224
rect -522 224 -518 228
rect -485 224 -481 228
rect -511 220 -507 224
rect -437 226 -433 230
rect -474 220 -470 224
rect -1382 138 -1377 143
rect -1898 106 -1894 110
rect -2176 88 -2172 92
rect -2166 84 -2162 88
rect -2144 88 -2140 92
rect -2107 88 -2103 92
rect -2133 84 -2129 88
rect -2059 90 -2055 94
rect -2096 84 -2092 88
rect -1865 107 -1861 111
rect -1832 99 -1827 104
rect -1818 91 -1813 96
rect -1781 91 -1777 95
rect -1746 99 -1741 104
rect -1368 130 -1363 135
rect -1353 121 -1348 126
rect -1320 125 -1316 129
rect -1012 126 -1008 130
rect -979 127 -975 131
rect -1732 91 -1727 96
rect -1695 91 -1691 95
rect -1665 94 -1661 98
rect -1654 94 -1650 98
rect -1627 93 -1623 97
rect -946 119 -941 124
rect -932 111 -927 116
rect -895 111 -891 115
rect -860 119 -855 124
rect -846 111 -841 116
rect -809 111 -805 115
rect -779 114 -775 118
rect -768 114 -764 118
rect -741 113 -737 117
rect -554 85 -550 89
rect -544 81 -540 85
rect -522 85 -518 89
rect -485 85 -481 89
rect -511 81 -507 85
rect -437 87 -433 91
rect -474 81 -470 85
rect -1700 11 -1695 16
rect -1686 3 -1681 8
rect -1649 3 -1645 7
rect -1378 18 -1373 23
rect -1364 10 -1359 15
rect -1327 10 -1323 14
rect -1290 18 -1286 22
rect -1279 18 -1275 22
rect -1252 17 -1248 21
rect -1012 9 -1008 13
rect -979 10 -975 14
rect -946 2 -941 7
rect -932 -6 -927 -1
rect -895 -6 -891 -2
rect -860 2 -855 7
rect -846 -6 -841 -1
rect -809 -6 -805 -2
rect -779 -3 -775 1
rect -768 -3 -764 1
rect -741 -4 -737 0
rect -562 -23 -558 -19
rect -552 -27 -548 -23
rect -530 -23 -526 -19
rect -493 -23 -489 -19
rect -519 -27 -515 -23
rect -445 -21 -441 -17
rect -482 -27 -478 -23
rect -2180 -58 -2176 -54
rect -2170 -62 -2166 -58
rect -2148 -58 -2144 -54
rect -2111 -58 -2107 -54
rect -2137 -62 -2133 -58
rect -2063 -56 -2059 -52
rect -2100 -62 -2096 -58
rect -2153 -186 -2149 -182
rect -2143 -190 -2139 -186
rect -2121 -186 -2117 -182
rect -2084 -186 -2080 -182
rect -2110 -190 -2106 -186
rect -2036 -184 -2032 -180
rect -2073 -190 -2069 -186
<< metal1 >>
rect -2164 836 -2041 840
rect -2158 830 -2154 836
rect -2126 825 -2122 836
rect -2090 825 -2086 836
rect -2048 832 -2023 836
rect -2041 826 -2037 832
rect -2138 791 -2134 810
rect -2103 802 -2099 815
rect -2067 804 -2063 815
rect -2033 804 -2029 816
rect -2103 798 -2088 802
rect -2067 800 -2040 804
rect -2033 800 -2021 804
rect -2103 791 -2099 798
rect -2067 791 -2063 800
rect -2033 797 -2029 800
rect -2158 775 -2154 786
rect -1906 793 -1881 797
rect -1873 794 -1848 798
rect -1838 797 -1769 801
rect -1752 797 -1683 801
rect -2041 783 -2037 792
rect -1899 787 -1895 793
rect -1866 788 -1862 794
rect -1838 789 -1833 797
rect -1807 789 -1802 797
rect -2126 775 -2122 781
rect -2090 775 -2086 781
rect -2045 779 -2025 783
rect -2045 775 -2041 779
rect -1775 782 -1770 797
rect -1752 789 -1747 797
rect -1721 789 -1716 797
rect -2158 769 -2041 775
rect -1891 765 -1887 777
rect -1858 766 -1854 778
rect -1906 761 -1898 765
rect -1891 761 -1879 765
rect -1873 762 -1865 766
rect -1858 762 -1846 766
rect -1891 758 -1887 761
rect -1858 759 -1854 762
rect -1824 759 -1819 779
rect -1789 778 -1764 782
rect -1689 782 -1684 797
rect -1672 788 -1623 792
rect -1666 782 -1662 788
rect -1629 784 -1623 788
rect -1782 772 -1778 778
rect -1835 754 -1832 759
rect -1824 755 -1802 759
rect -1899 744 -1895 753
rect -1866 745 -1862 754
rect -1835 746 -1818 751
rect -1807 750 -1802 755
rect -1774 750 -1770 762
rect -1738 759 -1733 779
rect -1703 778 -1678 782
rect -1696 772 -1692 778
rect -1632 780 -1610 784
rect -1628 774 -1624 780
rect -1749 754 -1746 759
rect -1738 755 -1716 759
rect -1807 746 -1781 750
rect -1774 746 -1762 750
rect -1749 746 -1732 751
rect -1721 750 -1716 755
rect -1688 750 -1684 762
rect -1721 746 -1695 750
rect -1688 746 -1676 750
rect -1647 752 -1643 762
rect -1620 752 -1616 764
rect -1647 748 -1627 752
rect -1620 748 -1608 752
rect -1903 740 -1883 744
rect -1870 741 -1850 745
rect -1807 742 -1802 746
rect -1774 743 -1770 746
rect -2162 735 -2039 739
rect -2156 729 -2152 735
rect -2124 724 -2120 735
rect -2088 724 -2084 735
rect -2046 731 -2021 735
rect -1721 742 -1716 746
rect -1688 743 -1684 746
rect -1647 745 -1643 748
rect -1620 745 -1616 748
rect -2039 725 -2035 731
rect -1838 728 -1833 732
rect -1782 729 -1778 738
rect -1657 742 -1643 745
rect -1657 738 -1653 742
rect -1786 728 -1766 729
rect -1838 725 -1766 728
rect -1752 728 -1747 732
rect -1696 729 -1692 738
rect -1700 728 -1680 729
rect -1752 725 -1680 728
rect -1666 727 -1662 733
rect -1647 731 -1643 733
rect -1628 731 -1624 740
rect -1647 727 -1612 731
rect -1838 724 -1802 725
rect -1752 724 -1716 725
rect -1666 724 -1643 727
rect -2136 690 -2132 709
rect -2101 701 -2097 714
rect -2065 703 -2061 714
rect -2031 703 -2027 715
rect -1706 709 -1637 713
rect -2101 697 -2086 701
rect -2065 699 -2038 703
rect -2031 699 -2019 703
rect -1706 701 -1701 709
rect -1675 701 -1670 709
rect -2101 690 -2097 697
rect -2065 690 -2061 699
rect -2031 696 -2027 699
rect -2156 674 -2152 685
rect -1643 694 -1638 709
rect -2039 682 -2035 691
rect -2124 674 -2120 680
rect -2088 674 -2084 680
rect -2043 678 -2023 682
rect -2043 674 -2039 678
rect -2156 668 -2039 674
rect -1692 671 -1687 691
rect -1657 690 -1632 694
rect -1650 684 -1646 690
rect -1703 666 -1700 671
rect -1692 667 -1670 671
rect -1703 658 -1686 663
rect -1675 662 -1670 667
rect -1642 662 -1638 674
rect -1675 658 -1649 662
rect -1642 658 -1630 662
rect -1675 654 -1670 658
rect -1642 655 -1638 658
rect -1706 640 -1701 644
rect -1650 641 -1646 650
rect -1654 640 -1634 641
rect -1706 637 -1634 640
rect -1363 639 -1294 643
rect -1706 636 -1670 637
rect -1363 631 -1358 639
rect -1332 631 -1327 639
rect -1300 624 -1295 639
rect -2175 610 -2052 614
rect -2169 604 -2165 610
rect -2137 599 -2133 610
rect -2101 599 -2097 610
rect -2059 606 -2034 610
rect -2052 600 -2048 606
rect -1349 601 -1344 621
rect -1314 620 -1289 624
rect -1307 614 -1303 620
rect -1360 596 -1357 601
rect -1349 597 -1327 601
rect -2149 565 -2145 584
rect -2114 576 -2110 589
rect -2078 578 -2074 589
rect -2044 578 -2040 590
rect -1908 581 -1883 585
rect -1875 582 -1850 586
rect -1840 585 -1771 589
rect -1754 585 -1685 589
rect -1360 588 -1343 593
rect -1332 592 -1327 597
rect -1299 592 -1295 604
rect -1332 588 -1306 592
rect -1299 588 -1266 592
rect -2114 572 -2099 576
rect -2078 574 -2051 578
rect -2044 574 -2032 578
rect -1901 575 -1897 581
rect -1868 576 -1864 582
rect -1840 577 -1835 585
rect -1809 577 -1804 585
rect -2114 565 -2110 572
rect -2078 565 -2074 574
rect -2044 571 -2040 574
rect -2169 549 -2165 560
rect -2052 557 -2048 566
rect -1777 570 -1772 585
rect -1754 577 -1749 585
rect -1723 577 -1718 585
rect -2137 549 -2133 555
rect -2101 549 -2097 555
rect -2056 553 -2036 557
rect -1893 553 -1889 565
rect -1860 554 -1856 566
rect -2056 549 -2052 553
rect -1908 549 -1900 553
rect -1893 549 -1881 553
rect -1875 550 -1867 554
rect -1860 550 -1848 554
rect -2169 543 -2052 549
rect -1893 546 -1889 549
rect -1860 547 -1856 550
rect -1826 547 -1821 567
rect -1791 566 -1766 570
rect -1691 570 -1686 585
rect -1332 584 -1327 588
rect -1299 585 -1295 588
rect -1674 576 -1625 580
rect -1668 570 -1664 576
rect -1631 572 -1625 576
rect -1784 560 -1780 566
rect -1837 542 -1834 547
rect -1826 543 -1804 547
rect -1901 532 -1897 541
rect -1868 533 -1864 542
rect -1837 534 -1820 539
rect -1809 538 -1804 543
rect -1776 538 -1772 550
rect -1740 547 -1735 567
rect -1705 566 -1680 570
rect -1698 560 -1694 566
rect -1634 568 -1612 572
rect -1363 570 -1358 574
rect -1307 571 -1303 580
rect -1311 570 -1291 571
rect -1630 562 -1626 568
rect -1363 567 -1291 570
rect -1363 566 -1327 567
rect -1751 542 -1748 547
rect -1740 543 -1718 547
rect -1809 534 -1783 538
rect -1776 534 -1764 538
rect -1751 534 -1734 539
rect -1723 538 -1718 543
rect -1690 538 -1686 550
rect -1723 534 -1697 538
rect -1690 534 -1678 538
rect -1649 540 -1645 550
rect -1622 540 -1618 552
rect -1649 536 -1629 540
rect -1622 536 -1610 540
rect -1367 538 -1295 542
rect -1905 528 -1885 532
rect -1872 529 -1852 533
rect -1809 530 -1804 534
rect -1776 531 -1772 534
rect -1723 530 -1718 534
rect -1690 531 -1686 534
rect -1649 533 -1645 536
rect -1622 533 -1618 536
rect -1840 516 -1835 520
rect -1784 517 -1780 526
rect -1659 530 -1645 533
rect -1659 526 -1655 530
rect -1367 530 -1362 538
rect -1336 530 -1331 538
rect -1788 516 -1768 517
rect -1840 513 -1768 516
rect -1754 516 -1749 520
rect -1698 517 -1694 526
rect -1702 516 -1682 517
rect -1754 513 -1682 516
rect -1668 515 -1664 521
rect -1649 519 -1645 521
rect -1630 519 -1626 528
rect -1301 522 -1296 538
rect -1649 515 -1614 519
rect -1840 512 -1804 513
rect -1754 512 -1718 513
rect -1668 512 -1645 515
rect -1708 497 -1639 501
rect -1353 500 -1348 520
rect -1324 500 -1320 520
rect -1310 518 -1285 522
rect -1708 489 -1703 497
rect -1677 489 -1672 497
rect -1645 482 -1640 497
rect -1353 496 -1320 500
rect -1303 508 -1299 518
rect -1324 486 -1320 496
rect -1295 486 -1291 498
rect -1269 500 -1266 588
rect -1234 554 -1165 558
rect -1234 548 -1230 554
rect -1172 538 -1165 554
rect -1172 534 -1150 538
rect -1168 528 -1164 534
rect -1269 496 -1233 500
rect -1194 499 -1188 508
rect -1160 506 -1156 518
rect -1175 502 -1167 506
rect -1160 502 -693 506
rect -1175 499 -1171 502
rect -1160 499 -1156 502
rect -1194 495 -1171 499
rect -1265 489 -1222 493
rect -1265 486 -1262 489
rect -2175 471 -2052 475
rect -2169 465 -2165 471
rect -2137 460 -2133 471
rect -2101 460 -2097 471
rect -2059 467 -2034 471
rect -2052 461 -2048 467
rect -1694 459 -1689 479
rect -1659 478 -1634 482
rect -1324 482 -1302 486
rect -1295 482 -1262 486
rect -1255 482 -1211 486
rect -1652 472 -1648 478
rect -1324 475 -1320 482
rect -1295 479 -1291 482
rect -1705 454 -1702 459
rect -1694 455 -1672 459
rect -2149 426 -2145 445
rect -2114 437 -2110 450
rect -2078 439 -2074 450
rect -2044 439 -2040 451
rect -1705 446 -1688 451
rect -1677 450 -1672 455
rect -1644 450 -1640 462
rect -1303 465 -1299 474
rect -1307 461 -1287 465
rect -1367 452 -1363 460
rect -1307 452 -1302 461
rect -1677 446 -1651 450
rect -1644 446 -1632 450
rect -1367 447 -1302 452
rect -1677 442 -1672 446
rect -1644 443 -1640 446
rect -2114 433 -2099 437
rect -2078 435 -2051 439
rect -2044 435 -2032 439
rect -2114 426 -2110 433
rect -2078 426 -2074 435
rect -2044 432 -2040 435
rect -2169 410 -2165 421
rect -1708 428 -1703 432
rect -1652 429 -1648 438
rect -1656 428 -1636 429
rect -2052 418 -2048 427
rect -1708 425 -1636 428
rect -1708 424 -1672 425
rect -2137 410 -2133 416
rect -2101 410 -2097 416
rect -2056 414 -2036 418
rect -1370 416 -1298 420
rect -2056 410 -2052 414
rect -2169 404 -2052 410
rect -1370 408 -1365 416
rect -1343 408 -1339 416
rect -1323 408 -1319 416
rect -1304 400 -1299 416
rect -1356 378 -1351 398
rect -1333 378 -1329 398
rect -1313 396 -1288 400
rect -1306 386 -1302 396
rect -2183 363 -2060 367
rect -1909 366 -1884 370
rect -1876 367 -1851 371
rect -1841 370 -1772 374
rect -1755 370 -1686 374
rect -1356 374 -1318 378
rect -2177 357 -2173 363
rect -2145 352 -2141 363
rect -2109 352 -2105 363
rect -2067 359 -2042 363
rect -1902 360 -1898 366
rect -1869 361 -1865 367
rect -1841 362 -1836 370
rect -1810 362 -1805 370
rect -2060 353 -2056 359
rect -1778 355 -1773 370
rect -1755 362 -1750 370
rect -1724 362 -1719 370
rect -2157 318 -2153 337
rect -2122 329 -2118 342
rect -2086 331 -2082 342
rect -2052 331 -2048 343
rect -1894 338 -1890 350
rect -1861 339 -1857 351
rect -1909 334 -1901 338
rect -1894 334 -1882 338
rect -1876 335 -1868 339
rect -1861 335 -1849 339
rect -1894 331 -1890 334
rect -1861 332 -1857 335
rect -1827 332 -1822 352
rect -1792 351 -1767 355
rect -1692 355 -1687 370
rect -1675 361 -1626 365
rect -1322 364 -1318 374
rect -1298 364 -1294 376
rect -1255 364 -1250 482
rect -1194 479 -1188 495
rect -1224 476 -1188 479
rect -1224 473 -1220 476
rect -1203 473 -1199 476
rect -1234 464 -1230 468
rect -1212 464 -1208 468
rect -1194 464 -1188 468
rect -1168 464 -1164 494
rect -1234 461 -1164 464
rect -696 454 -693 502
rect -550 488 -427 492
rect -544 482 -540 488
rect -512 477 -508 488
rect -476 477 -472 488
rect -434 484 -409 488
rect -427 478 -423 484
rect -696 450 -543 454
rect -524 443 -520 462
rect -489 454 -485 467
rect -453 456 -449 467
rect -419 456 -415 468
rect -489 450 -474 454
rect -453 452 -426 456
rect -419 452 -407 456
rect -489 443 -485 450
rect -453 443 -449 452
rect -419 449 -415 452
rect -544 427 -540 438
rect -427 435 -423 444
rect -512 427 -508 433
rect -476 427 -472 433
rect -431 431 -411 435
rect -431 427 -427 431
rect -544 421 -427 427
rect -1018 395 -993 399
rect -985 396 -960 400
rect -950 399 -881 403
rect -864 399 -795 403
rect -1011 389 -1007 395
rect -978 390 -974 396
rect -950 391 -945 399
rect -919 391 -914 399
rect -887 384 -882 399
rect -864 391 -859 399
rect -833 391 -828 399
rect -1003 367 -999 379
rect -970 368 -966 380
rect -1669 355 -1665 361
rect -1632 357 -1626 361
rect -1322 360 -1305 364
rect -1298 360 -1250 364
rect -1018 363 -1010 367
rect -1003 363 -991 367
rect -985 364 -977 368
rect -970 364 -958 368
rect -1003 360 -999 363
rect -970 361 -966 364
rect -936 361 -931 381
rect -901 380 -876 384
rect -801 384 -796 399
rect -784 390 -735 394
rect -778 384 -774 390
rect -741 386 -735 390
rect -548 387 -425 391
rect -894 374 -890 380
rect -1785 345 -1781 351
rect -2122 325 -2107 329
rect -2086 327 -2059 331
rect -2052 327 -2040 331
rect -2122 318 -2118 325
rect -2086 318 -2082 327
rect -2052 324 -2048 327
rect -2177 302 -2173 313
rect -1838 327 -1835 332
rect -1827 328 -1805 332
rect -2060 310 -2056 319
rect -1902 317 -1898 326
rect -1869 318 -1865 327
rect -1838 319 -1821 324
rect -1810 323 -1805 328
rect -1777 323 -1773 335
rect -1741 332 -1736 352
rect -1706 351 -1681 355
rect -1699 345 -1695 351
rect -1635 353 -1613 357
rect -1322 353 -1318 360
rect -1298 357 -1294 360
rect -1631 347 -1627 353
rect -1752 327 -1749 332
rect -1741 328 -1719 332
rect -1810 319 -1784 323
rect -1777 319 -1765 323
rect -1752 319 -1735 324
rect -1724 323 -1719 328
rect -1691 323 -1687 335
rect -1724 319 -1698 323
rect -1691 319 -1679 323
rect -1650 325 -1646 335
rect -1623 325 -1619 337
rect -947 356 -944 361
rect -936 357 -914 361
rect -1306 343 -1302 352
rect -1011 346 -1007 355
rect -978 347 -974 356
rect -947 348 -930 353
rect -919 352 -914 357
rect -886 352 -882 364
rect -850 361 -845 381
rect -815 380 -790 384
rect -808 374 -804 380
rect -744 382 -722 386
rect -740 376 -736 382
rect -542 381 -538 387
rect -861 356 -858 361
rect -850 357 -828 361
rect -919 348 -893 352
rect -886 348 -874 352
rect -861 348 -844 353
rect -833 352 -828 357
rect -800 352 -796 364
rect -833 348 -807 352
rect -800 348 -788 352
rect -759 354 -755 364
rect -732 354 -728 366
rect -510 376 -506 387
rect -474 376 -470 387
rect -432 383 -407 387
rect -425 377 -421 383
rect -759 350 -739 354
rect -732 353 -572 354
rect -732 350 -541 353
rect -1310 339 -1290 343
rect -1015 342 -995 346
rect -982 343 -962 347
rect -919 344 -914 348
rect -886 345 -882 348
rect -1370 329 -1366 333
rect -1310 329 -1305 339
rect -1370 325 -1305 329
rect -833 344 -828 348
rect -800 345 -796 348
rect -759 347 -755 350
rect -732 347 -728 350
rect -575 349 -541 350
rect -950 330 -945 334
rect -894 331 -890 340
rect -769 344 -755 347
rect -769 340 -765 344
rect -522 342 -518 361
rect -487 353 -483 366
rect -451 355 -447 366
rect -417 355 -413 367
rect -487 349 -472 353
rect -451 351 -424 355
rect -417 351 -405 355
rect -487 342 -483 349
rect -451 342 -447 351
rect -417 348 -413 351
rect -898 330 -878 331
rect -950 327 -878 330
rect -864 330 -859 334
rect -808 331 -804 340
rect -812 330 -792 331
rect -864 327 -792 330
rect -778 329 -774 335
rect -759 333 -755 335
rect -740 333 -736 342
rect -759 329 -724 333
rect -950 326 -914 327
rect -864 326 -828 327
rect -778 326 -755 329
rect -542 326 -538 337
rect -425 334 -421 343
rect -510 326 -506 332
rect -474 326 -470 332
rect -429 330 -409 334
rect -429 326 -425 330
rect -1650 321 -1630 325
rect -1623 321 -1611 325
rect -1906 313 -1886 317
rect -1873 314 -1853 318
rect -1810 315 -1805 319
rect -1777 316 -1773 319
rect -2145 302 -2141 308
rect -2109 302 -2105 308
rect -2064 306 -2044 310
rect -2064 302 -2060 306
rect -2177 296 -2060 302
rect -1724 315 -1719 319
rect -1691 316 -1687 319
rect -1650 318 -1646 321
rect -1623 318 -1619 321
rect -542 320 -425 326
rect -1841 301 -1836 305
rect -1785 302 -1781 311
rect -1660 315 -1646 318
rect -1660 311 -1656 315
rect -1789 301 -1769 302
rect -1841 298 -1769 301
rect -1755 301 -1750 305
rect -1699 302 -1695 311
rect -1703 301 -1683 302
rect -1755 298 -1683 301
rect -1669 300 -1665 306
rect -1650 304 -1646 306
rect -1631 304 -1627 313
rect -1650 300 -1615 304
rect -1841 297 -1805 298
rect -1755 297 -1719 298
rect -1669 297 -1646 300
rect -1709 282 -1640 286
rect -1381 282 -1312 286
rect -1709 274 -1704 282
rect -1678 274 -1673 282
rect -1646 267 -1641 282
rect -1381 274 -1376 282
rect -1350 274 -1345 282
rect -2189 254 -2066 258
rect -2183 248 -2179 254
rect -2151 243 -2147 254
rect -2115 243 -2111 254
rect -2073 250 -2048 254
rect -2066 244 -2062 250
rect -1695 244 -1690 264
rect -1660 263 -1635 267
rect -1318 267 -1313 282
rect -1018 278 -993 282
rect -985 279 -960 283
rect -950 282 -881 286
rect -864 282 -795 286
rect -1011 272 -1007 278
rect -978 273 -974 279
rect -950 274 -945 282
rect -919 274 -914 282
rect -1653 257 -1649 263
rect -1706 239 -1703 244
rect -1695 240 -1673 244
rect -2163 209 -2159 228
rect -2128 220 -2124 233
rect -2092 222 -2088 233
rect -2058 222 -2054 234
rect -1706 231 -1689 236
rect -1678 235 -1673 240
rect -1645 235 -1641 247
rect -1367 244 -1362 264
rect -1332 263 -1307 267
rect -1325 257 -1321 263
rect -887 267 -882 282
rect -864 274 -859 282
rect -833 274 -828 282
rect -1279 253 -1203 257
rect -1378 239 -1375 244
rect -1367 240 -1345 244
rect -1678 231 -1652 235
rect -1645 231 -1633 235
rect -1378 231 -1361 236
rect -1350 235 -1345 240
rect -1317 235 -1313 247
rect -1273 245 -1269 253
rect -1350 231 -1324 235
rect -1317 231 -1298 235
rect -1678 227 -1673 231
rect -1645 228 -1641 231
rect -2128 216 -2113 220
rect -2092 218 -2065 222
rect -2058 218 -2046 222
rect -2128 209 -2124 216
rect -2092 209 -2088 218
rect -2058 215 -2054 218
rect -2183 193 -2179 204
rect -1350 227 -1345 231
rect -1317 228 -1313 231
rect -1709 213 -1704 217
rect -1653 214 -1649 223
rect -1657 213 -1637 214
rect -1709 210 -1637 213
rect -1381 213 -1376 217
rect -1325 214 -1321 223
rect -1329 213 -1309 214
rect -1381 210 -1309 213
rect -2066 201 -2062 210
rect -1709 209 -1673 210
rect -1381 209 -1345 210
rect -1302 206 -1298 231
rect -1211 244 -1204 253
rect -1003 250 -999 262
rect -970 251 -966 263
rect -1018 246 -1010 250
rect -1003 246 -991 250
rect -985 247 -977 251
rect -970 247 -958 251
rect -1211 240 -1189 244
rect -1003 243 -999 246
rect -970 244 -966 247
rect -936 244 -931 264
rect -901 263 -876 267
rect -801 267 -796 282
rect -784 273 -735 277
rect -778 267 -774 273
rect -741 269 -735 273
rect -894 257 -890 263
rect -1207 234 -1203 240
rect -947 239 -944 244
rect -936 240 -914 244
rect -1011 229 -1007 238
rect -978 230 -974 239
rect -947 231 -930 236
rect -919 235 -914 240
rect -886 235 -882 247
rect -850 244 -845 264
rect -815 263 -790 267
rect -808 257 -804 263
rect -744 265 -722 269
rect -740 259 -736 265
rect -561 262 -438 266
rect -861 239 -858 244
rect -850 240 -828 244
rect -919 231 -893 235
rect -886 231 -874 235
rect -861 231 -844 236
rect -833 235 -828 240
rect -800 235 -796 247
rect -833 231 -807 235
rect -800 231 -788 235
rect -759 237 -755 247
rect -732 237 -728 249
rect -555 256 -551 262
rect -759 233 -739 237
rect -732 233 -598 237
rect -523 251 -519 262
rect -487 251 -483 262
rect -445 258 -420 262
rect -438 252 -434 258
rect -1015 225 -995 229
rect -982 226 -962 230
rect -919 227 -914 231
rect -886 228 -882 231
rect -1302 202 -1272 206
rect -1233 205 -1227 215
rect -1199 212 -1195 224
rect -833 227 -828 231
rect -800 228 -796 231
rect -759 230 -755 233
rect -732 230 -728 233
rect -950 213 -945 217
rect -894 214 -890 223
rect -769 227 -755 230
rect -769 223 -765 227
rect -601 228 -598 233
rect -898 213 -878 214
rect -1214 208 -1206 212
rect -1199 208 -1187 212
rect -950 210 -878 213
rect -864 213 -859 217
rect -808 214 -804 223
rect -812 213 -792 214
rect -864 210 -792 213
rect -778 212 -774 218
rect -759 216 -755 218
rect -740 216 -736 225
rect -601 224 -554 228
rect -535 217 -531 236
rect -500 228 -496 241
rect -464 230 -460 241
rect -430 230 -426 242
rect -500 224 -485 228
rect -464 226 -437 230
rect -430 226 -418 230
rect -500 217 -496 224
rect -464 217 -460 226
rect -430 223 -426 226
rect -759 212 -724 216
rect -950 209 -914 210
rect -864 209 -828 210
rect -778 209 -755 212
rect -1214 205 -1210 208
rect -1199 205 -1195 208
rect -1233 201 -1210 205
rect -2151 193 -2147 199
rect -2115 193 -2111 199
rect -2070 197 -2050 201
rect -2070 193 -2066 197
rect -2183 187 -2066 193
rect -1285 189 -1248 193
rect -1385 181 -1313 185
rect -1385 173 -1380 181
rect -1354 173 -1349 181
rect -1319 165 -1314 181
rect -1906 138 -1881 142
rect -1873 139 -1848 143
rect -1838 142 -1769 146
rect -1752 142 -1683 146
rect -1371 143 -1366 163
rect -1342 143 -1338 163
rect -1328 161 -1303 165
rect -1899 132 -1895 138
rect -1866 133 -1862 139
rect -1838 134 -1833 142
rect -1807 134 -1802 142
rect -2183 126 -2060 130
rect -2177 120 -2173 126
rect -2145 115 -2141 126
rect -2109 115 -2105 126
rect -2067 122 -2042 126
rect -1775 127 -1770 142
rect -1752 134 -1747 142
rect -1721 134 -1716 142
rect -2060 116 -2056 122
rect -1891 110 -1887 122
rect -1858 111 -1854 123
rect -1906 106 -1898 110
rect -1891 106 -1879 110
rect -1873 107 -1865 111
rect -1858 107 -1846 111
rect -2157 81 -2153 100
rect -2122 92 -2118 105
rect -2086 94 -2082 105
rect -2052 94 -2048 106
rect -1891 103 -1887 106
rect -1858 104 -1854 107
rect -1824 104 -1819 124
rect -1789 123 -1764 127
rect -1689 127 -1684 142
rect -1371 139 -1338 143
rect -1321 151 -1317 161
rect -1672 133 -1623 137
rect -1666 127 -1662 133
rect -1629 129 -1623 133
rect -1342 129 -1338 139
rect -1313 129 -1309 141
rect -1285 129 -1282 189
rect -1233 186 -1227 201
rect -1263 183 -1227 186
rect -1263 180 -1259 183
rect -1233 180 -1227 183
rect -555 201 -551 212
rect -438 209 -434 218
rect -523 201 -519 207
rect -487 201 -483 207
rect -442 205 -422 209
rect -442 201 -438 205
rect -1273 170 -1269 176
rect -1251 170 -1247 176
rect -1207 170 -1203 200
rect -555 195 -438 201
rect -1273 167 -1203 170
rect -1020 158 -995 162
rect -987 159 -962 163
rect -952 162 -883 166
rect -866 162 -797 166
rect -1013 152 -1009 158
rect -980 153 -976 159
rect -952 154 -947 162
rect -921 154 -916 162
rect -889 147 -884 162
rect -866 154 -861 162
rect -835 154 -830 162
rect -1005 130 -1001 142
rect -972 131 -968 143
rect -1782 117 -1778 123
rect -1835 99 -1832 104
rect -1824 100 -1802 104
rect -2122 88 -2107 92
rect -2086 90 -2059 94
rect -2052 90 -2040 94
rect -2122 81 -2118 88
rect -2086 81 -2082 90
rect -2052 87 -2048 90
rect -1899 89 -1895 98
rect -1866 90 -1862 99
rect -1835 91 -1818 96
rect -1807 95 -1802 100
rect -1774 95 -1770 107
rect -1738 104 -1733 124
rect -1703 123 -1678 127
rect -1696 117 -1692 123
rect -1632 125 -1610 129
rect -1628 119 -1624 125
rect -1425 121 -1353 126
rect -1342 125 -1320 129
rect -1313 125 -1282 129
rect -1020 126 -1012 130
rect -1005 126 -993 130
rect -987 127 -979 131
rect -972 127 -960 131
rect -1749 99 -1746 104
rect -1738 100 -1716 104
rect -1807 91 -1781 95
rect -1774 91 -1762 95
rect -1749 91 -1732 96
rect -1721 95 -1716 100
rect -1688 95 -1684 107
rect -1721 91 -1695 95
rect -1688 91 -1676 95
rect -1647 97 -1643 107
rect -1620 97 -1616 109
rect -1647 93 -1627 97
rect -1620 93 -1608 97
rect -2177 65 -2173 76
rect -1903 85 -1883 89
rect -1870 86 -1850 90
rect -1807 87 -1802 91
rect -1774 88 -1770 91
rect -2060 73 -2056 82
rect -1721 87 -1716 91
rect -1688 88 -1684 91
rect -1647 90 -1643 93
rect -1620 90 -1616 93
rect -1838 73 -1833 77
rect -1782 74 -1778 83
rect -1657 87 -1643 90
rect -1657 83 -1653 87
rect -1786 73 -1766 74
rect -2145 65 -2141 71
rect -2109 65 -2105 71
rect -2064 69 -2044 73
rect -1838 70 -1766 73
rect -1752 73 -1747 77
rect -1696 74 -1692 83
rect -1700 73 -1680 74
rect -1752 70 -1680 73
rect -1666 72 -1662 78
rect -1647 76 -1643 78
rect -1628 76 -1624 85
rect -1647 72 -1612 76
rect -1838 69 -1802 70
rect -1752 69 -1716 70
rect -1666 69 -1643 72
rect -2064 65 -2060 69
rect -2177 59 -2060 65
rect -1706 54 -1637 58
rect -1706 46 -1701 54
rect -1675 46 -1670 54
rect -1643 39 -1638 54
rect -1692 16 -1687 36
rect -1657 35 -1632 39
rect -1650 29 -1646 35
rect -1703 11 -1700 16
rect -1692 12 -1670 16
rect -1703 3 -1686 8
rect -1675 7 -1670 12
rect -1642 7 -1638 19
rect -1425 7 -1419 121
rect -1342 118 -1338 125
rect -1313 122 -1309 125
rect -1005 123 -1001 126
rect -972 124 -968 127
rect -938 124 -933 144
rect -903 143 -878 147
rect -803 147 -798 162
rect -786 153 -737 157
rect -780 147 -776 153
rect -743 149 -737 153
rect -896 137 -892 143
rect -949 119 -946 124
rect -938 120 -916 124
rect -1321 108 -1317 117
rect -1013 109 -1009 118
rect -980 110 -976 119
rect -949 111 -932 116
rect -921 115 -916 120
rect -888 115 -884 127
rect -852 124 -847 144
rect -817 143 -792 147
rect -810 137 -806 143
rect -746 145 -724 149
rect -742 139 -738 145
rect -863 119 -860 124
rect -852 120 -830 124
rect -921 111 -895 115
rect -888 111 -876 115
rect -863 111 -846 116
rect -835 115 -830 120
rect -802 115 -798 127
rect -835 111 -809 115
rect -802 111 -790 115
rect -761 117 -757 127
rect -734 117 -730 129
rect -561 123 -438 127
rect -555 117 -551 123
rect -761 113 -741 117
rect -734 113 -596 117
rect -1325 104 -1305 108
rect -1017 105 -997 109
rect -984 106 -964 110
rect -921 107 -916 111
rect -888 108 -884 111
rect -1385 95 -1381 103
rect -1325 95 -1320 104
rect -1385 90 -1320 95
rect -835 107 -830 111
rect -802 108 -798 111
rect -761 110 -757 113
rect -734 110 -730 113
rect -952 93 -947 97
rect -896 94 -892 103
rect -771 107 -757 110
rect -771 103 -767 107
rect -900 93 -880 94
rect -952 90 -880 93
rect -866 93 -861 97
rect -810 94 -806 103
rect -814 93 -794 94
rect -866 90 -794 93
rect -780 92 -776 98
rect -761 96 -757 98
rect -742 96 -738 105
rect -761 92 -726 96
rect -952 89 -916 90
rect -866 89 -830 90
rect -780 89 -757 92
rect -600 89 -596 113
rect -523 112 -519 123
rect -487 112 -483 123
rect -445 119 -420 123
rect -438 113 -434 119
rect -600 85 -554 89
rect -535 78 -531 97
rect -500 89 -496 102
rect -464 91 -460 102
rect -430 91 -426 103
rect -500 85 -485 89
rect -464 87 -437 91
rect -430 87 -418 91
rect -500 78 -496 85
rect -464 78 -460 87
rect -430 84 -426 87
rect -1384 61 -1315 65
rect -555 62 -551 73
rect -438 70 -434 79
rect -523 62 -519 68
rect -487 62 -483 68
rect -442 66 -422 70
rect -442 62 -438 66
rect -1384 53 -1379 61
rect -1353 53 -1348 61
rect -1321 46 -1316 61
rect -1297 57 -1248 61
rect -1291 51 -1287 57
rect -1254 53 -1248 57
rect -555 56 -438 62
rect -1370 23 -1365 43
rect -1335 42 -1310 46
rect -1328 36 -1324 42
rect -1257 49 -1235 53
rect -1253 43 -1249 49
rect -1020 41 -995 45
rect -987 42 -962 46
rect -952 45 -883 49
rect -866 45 -797 49
rect -1381 18 -1378 23
rect -1370 19 -1348 23
rect -1381 13 -1364 15
rect -1406 10 -1364 13
rect -1353 14 -1348 19
rect -1320 14 -1316 26
rect -1302 18 -1290 22
rect -1272 21 -1268 31
rect -1245 21 -1241 33
rect -1013 35 -1009 41
rect -980 36 -976 42
rect -952 37 -947 45
rect -921 37 -916 45
rect -889 30 -884 45
rect -866 37 -861 45
rect -835 37 -830 45
rect -1302 14 -1299 18
rect -1272 17 -1252 21
rect -1245 17 -1233 21
rect -1272 14 -1268 17
rect -1245 14 -1241 17
rect -1353 10 -1327 14
rect -1320 10 -1299 14
rect -1282 11 -1268 14
rect -1406 7 -1403 10
rect -1675 3 -1649 7
rect -1642 3 -1403 7
rect -1353 6 -1348 10
rect -1320 7 -1316 10
rect -1282 7 -1278 11
rect -1005 13 -1001 25
rect -972 14 -968 26
rect -1020 9 -1012 13
rect -1005 9 -993 13
rect -987 10 -979 14
rect -972 10 -960 14
rect -1675 -1 -1670 3
rect -1642 0 -1638 3
rect -1706 -15 -1701 -11
rect -1650 -14 -1646 -5
rect -1384 -8 -1379 -4
rect -1328 -7 -1324 2
rect -1291 -4 -1287 2
rect -1272 0 -1268 2
rect -1253 0 -1249 9
rect -1005 6 -1001 9
rect -972 7 -968 10
rect -938 7 -933 27
rect -903 26 -878 30
rect -803 30 -798 45
rect -786 36 -737 40
rect -780 30 -776 36
rect -743 32 -737 36
rect -896 20 -892 26
rect -949 2 -946 7
rect -938 3 -916 7
rect -1272 -4 -1237 0
rect -1291 -7 -1268 -4
rect -1332 -8 -1312 -7
rect -1013 -8 -1009 1
rect -980 -7 -976 2
rect -949 -6 -932 -1
rect -921 -2 -916 3
rect -888 -2 -884 10
rect -852 7 -847 27
rect -817 26 -792 30
rect -810 20 -806 26
rect -746 28 -724 32
rect -742 22 -738 28
rect -569 15 -446 19
rect -863 2 -860 7
rect -852 3 -830 7
rect -921 -6 -895 -2
rect -888 -6 -876 -2
rect -863 -6 -846 -1
rect -835 -2 -830 3
rect -802 -2 -798 10
rect -835 -6 -809 -2
rect -802 -6 -790 -2
rect -761 0 -757 10
rect -734 0 -730 12
rect -563 9 -559 15
rect -761 -4 -741 0
rect -734 -4 -613 0
rect -1384 -11 -1312 -8
rect -1384 -12 -1348 -11
rect -1017 -12 -997 -8
rect -984 -11 -964 -7
rect -921 -10 -916 -6
rect -888 -9 -884 -6
rect -1654 -15 -1634 -14
rect -2187 -20 -2064 -16
rect -1706 -18 -1634 -15
rect -1706 -19 -1670 -18
rect -835 -10 -830 -6
rect -802 -9 -798 -6
rect -761 -7 -757 -4
rect -734 -7 -730 -4
rect -2181 -26 -2177 -20
rect -2149 -31 -2145 -20
rect -2113 -31 -2109 -20
rect -2071 -24 -2046 -20
rect -952 -24 -947 -20
rect -896 -23 -892 -14
rect -771 -10 -757 -7
rect -771 -14 -767 -10
rect -900 -24 -880 -23
rect -2064 -30 -2060 -24
rect -952 -27 -880 -24
rect -866 -24 -861 -20
rect -810 -23 -806 -14
rect -814 -24 -794 -23
rect -866 -27 -794 -24
rect -780 -25 -776 -19
rect -761 -21 -757 -19
rect -742 -21 -738 -12
rect -616 -19 -613 -4
rect -531 4 -527 15
rect -495 4 -491 15
rect -453 11 -428 15
rect -446 5 -442 11
rect -761 -25 -726 -21
rect -616 -23 -562 -19
rect -952 -28 -916 -27
rect -866 -28 -830 -27
rect -780 -28 -757 -25
rect -543 -30 -539 -11
rect -508 -19 -504 -6
rect -472 -17 -468 -6
rect -438 -17 -434 -5
rect -508 -23 -493 -19
rect -472 -21 -445 -17
rect -438 -21 -426 -17
rect -508 -30 -504 -23
rect -472 -30 -468 -21
rect -438 -24 -434 -21
rect -2161 -65 -2157 -46
rect -2126 -54 -2122 -41
rect -2090 -52 -2086 -41
rect -2056 -52 -2052 -40
rect -563 -46 -559 -35
rect -446 -38 -442 -29
rect -531 -46 -527 -40
rect -495 -46 -491 -40
rect -450 -42 -430 -38
rect -450 -46 -446 -42
rect -563 -52 -446 -46
rect -2126 -58 -2111 -54
rect -2090 -56 -2063 -52
rect -2056 -56 -2044 -52
rect -2126 -65 -2122 -58
rect -2090 -65 -2086 -56
rect -2056 -59 -2052 -56
rect -2181 -81 -2177 -70
rect -2064 -73 -2060 -64
rect -2149 -81 -2145 -75
rect -2113 -81 -2109 -75
rect -2068 -77 -2048 -73
rect -2068 -81 -2064 -77
rect -2181 -87 -2064 -81
rect -2160 -148 -2037 -144
rect -2154 -154 -2150 -148
rect -2122 -159 -2118 -148
rect -2086 -159 -2082 -148
rect -2044 -152 -2019 -148
rect -2037 -158 -2033 -152
rect -2134 -193 -2130 -174
rect -2099 -182 -2095 -169
rect -2063 -180 -2059 -169
rect -2029 -180 -2025 -168
rect -2099 -186 -2084 -182
rect -2063 -184 -2036 -180
rect -2029 -184 -2017 -180
rect -2099 -193 -2095 -186
rect -2063 -193 -2059 -184
rect -2029 -187 -2025 -184
rect -2154 -209 -2150 -198
rect -2037 -201 -2033 -192
rect -2122 -209 -2118 -203
rect -2086 -209 -2082 -203
rect -2041 -205 -2021 -201
rect -2041 -209 -2037 -205
rect -2154 -215 -2037 -209
<< labels >>
rlabel pdcontact -1326 31 -1326 31 1 vdd
rlabel ndcontact -1326 4 -1326 4 1 gnd
rlabel metal1 -1324 -9 -1324 -9 1 gnd
rlabel metal1 -1368 63 -1368 63 5 vdd
rlabel ndcontact -1382 4 -1382 4 1 gnd
rlabel pdcontact -1382 48 -1382 48 1 vdd
rlabel pdcontact -1351 47 -1351 47 1 vdd
rlabel polycontact -1375 20 -1375 20 1 p1
rlabel polycontact -1361 12 -1361 12 1 g0
rlabel ndiffusion -1368 1 -1368 1 1 n29
rlabel metal1 -1311 12 -1311 12 7 p1g0
rlabel ndcontact -1318 4 -1318 4 1 p1g0
rlabel pdcontact -1318 31 -1318 31 1 p1g0
rlabel polycontact -1325 12 -1325 12 1 nand17
rlabel ndcontact -1351 1 -1351 1 1 nand17
rlabel pdcontact -1368 48 -1368 48 1 nand17
rlabel pdcontact -1251 38 -1251 38 1 vdd
rlabel ndcontact -1251 11 -1251 11 1 gnd
rlabel metal1 -1280 -6 -1280 -6 1 gnd
rlabel metal1 -1280 59 -1280 59 5 vdd
rlabel pdcontact -1289 41 -1289 41 1 vdd
rlabel ndcontact -1271 4 -1271 4 1 gnd
rlabel ndcontact -1289 5 -1289 5 1 gnd
rlabel polycontact -1250 19 -1250 19 1 nor9
rlabel pdcontact -1270 41 -1270 41 1 nor9
rlabel ndcontact -1280 4 -1280 4 1 nor9
rlabel pdiffusion -1280 42 -1280 42 1 n30
rlabel polycontact -1288 20 -1288 20 1 p1g0
rlabel polycontact -1277 20 -1277 20 1 g1
rlabel metal1 -1236 19 -1236 19 7 c2
rlabel ndcontact -1243 11 -1243 11 1 c2
rlabel pdcontact -1243 38 -1243 38 1 c2
rlabel metal1 -1369 183 -1369 183 5 vdd
rlabel pdcontact -1383 168 -1383 168 1 vdd
rlabel pdcontact -1352 168 -1352 168 1 vdd
rlabel ndcontact -1383 110 -1383 110 1 gnd
rlabel pdcontact -1319 146 -1319 146 1 vdd
rlabel ndcontact -1319 119 -1319 119 1 gnd
rlabel metal1 -1317 106 -1317 106 1 gnd
rlabel pdcontact -1323 252 -1323 252 1 vdd
rlabel ndcontact -1323 225 -1323 225 1 gnd
rlabel metal1 -1321 212 -1321 212 1 gnd
rlabel metal1 -1365 284 -1365 284 5 vdd
rlabel ndcontact -1379 225 -1379 225 1 gnd
rlabel pdcontact -1379 269 -1379 269 1 vdd
rlabel pdcontact -1348 268 -1348 268 1 vdd
rlabel metal1 -1257 255 -1257 255 5 vdd
rlabel pdcontact -1271 230 -1271 230 1 vdd
rlabel pdcontact -1205 229 -1205 229 1 vdd
rlabel ndcontact -1205 202 -1205 202 1 gnd
rlabel ndcontact -1271 178 -1271 178 1 gnd
rlabel ndcontact -1249 178 -1249 178 1 gnd
rlabel metal1 -1236 168 -1236 168 1 gnd
rlabel metal1 -1354 418 -1354 418 5 vdd
rlabel pdcontact -1368 403 -1368 403 1 vdd
rlabel ndcontact -1368 345 -1368 345 1 gnd
rlabel pdcontact -1304 381 -1304 381 1 vdd
rlabel ndcontact -1304 354 -1304 354 1 gnd
rlabel metal1 -1302 341 -1302 341 1 gnd
rlabel pdcontact -1341 402 -1341 402 1 vdd
rlabel pdcontact -1321 403 -1321 403 1 vdd
rlabel metal1 -1351 540 -1351 540 5 vdd
rlabel pdcontact -1365 525 -1365 525 1 vdd
rlabel pdcontact -1334 525 -1334 525 1 vdd
rlabel ndcontact -1365 467 -1365 467 1 gnd
rlabel pdcontact -1301 503 -1301 503 1 vdd
rlabel ndcontact -1301 476 -1301 476 1 gnd
rlabel metal1 -1299 463 -1299 463 1 gnd
rlabel pdcontact -1305 609 -1305 609 1 vdd
rlabel ndcontact -1305 582 -1305 582 1 gnd
rlabel metal1 -1303 569 -1303 569 1 gnd
rlabel metal1 -1347 641 -1347 641 5 vdd
rlabel ndcontact -1361 582 -1361 582 1 gnd
rlabel pdcontact -1361 626 -1361 626 1 vdd
rlabel pdcontact -1330 625 -1330 625 1 vdd
rlabel pdcontact -1232 524 -1232 524 1 vdd
rlabel pdcontact -1166 523 -1166 523 1 vdd
rlabel ndcontact -1166 496 -1166 496 1 gnd
rlabel ndcontact -1232 472 -1232 472 1 gnd
rlabel ndcontact -1210 472 -1210 472 1 gnd
rlabel metal1 -1197 462 -1197 462 1 gnd
rlabel ndcontact -1191 472 -1191 472 1 gnd
rlabel metal1 -1190 556 -1190 556 5 vdd
rlabel polycontact -1379 140 -1379 140 1 p2
rlabel polycontact -1366 132 -1366 132 1 p1
rlabel polycontact -1350 124 -1350 124 1 g0
rlabel ndiffusion -1368 111 -1368 111 1 n31
rlabel ndiffusion -1353 111 -1353 111 1 n32
rlabel ndcontact -1340 110 -1340 110 1 nand18
rlabel polycontact -1318 127 -1318 127 1 nand18
rlabel pdcontact -1340 168 -1340 168 1 nand18
rlabel pdcontact -1369 167 -1369 167 1 nand18
rlabel metal1 -1304 127 -1304 127 1 p2p1g0
rlabel pdcontact -1311 146 -1311 146 1 p2p1g0
rlabel ndcontact -1311 119 -1311 119 1 p2p1g0
rlabel polycontact -1372 241 -1372 241 1 p2
rlabel polycontact -1358 233 -1358 233 1 g1
rlabel ndiffusion -1365 222 -1365 222 1 n33
rlabel polycontact -1322 233 -1322 233 1 nand19
rlabel ndcontact -1348 222 -1348 222 1 nand19
rlabel pdcontact -1365 269 -1365 269 1 nand19
rlabel metal1 -1309 233 -1309 233 1 p2g1
rlabel pdcontact -1315 252 -1315 252 1 p2g1
rlabel ndcontact -1315 225 -1315 225 1 p2g1
rlabel polycontact -1270 204 -1270 204 1 p2g1
rlabel polycontact -1246 191 -1246 191 1 p2p1g0
rlabel polycontact -1259 198 -1259 198 1 g2
rlabel metal1 -1190 210 -1190 210 1 c3
rlabel pdcontact -1197 229 -1197 229 1 c3
rlabel ndcontact -1197 202 -1197 202 1 c3
rlabel pdiffusion -1262 230 -1262 230 1 n34
rlabel pdiffusion -1250 229 -1250 229 1 n35
rlabel polycontact -1204 210 -1204 210 1 nor10
rlabel pdcontact -1230 230 -1230 230 1 nor10
rlabel ndcontact -1230 178 -1230 178 1 nor10
rlabel polycontact -1165 504 -1165 504 1 nor11
rlabel pdcontact -1191 524 -1191 524 1 nor11
rlabel ndcontact -1261 178 -1261 178 1 nor10
rlabel ndcontact -1201 472 -1201 472 1 nor11
rlabel ndcontact -1222 472 -1222 472 1 nor11
rlabel metal1 -1151 504 -1151 504 7 c4
rlabel ndcontact -1158 496 -1158 496 1 c4
rlabel pdcontact -1158 523 -1158 523 1 c4
rlabel ndiffusion -1353 346 -1353 346 1 n36
rlabel ndiffusion -1338 346 -1338 346 1 n37
rlabel ndiffusion -1331 345 -1331 345 1 n38
rlabel ndiffusion -1350 468 -1350 468 1 n39
rlabel ndiffusion -1335 468 -1335 468 1 n40
rlabel ndiffusion -1347 579 -1347 579 1 n41
rlabel pdiffusion -1223 524 -1223 524 1 n42
rlabel pdiffusion -1211 523 -1211 523 1 n43
rlabel pdiffusion -1201 524 -1201 524 1 n44
rlabel polycontact -1303 362 -1303 362 1 nand20
rlabel ndcontact -1320 342 -1320 342 1 nand20
rlabel pdcontact -1331 403 -1331 403 1 nand20
rlabel pdcontact -1354 402 -1354 402 1 nand20
rlabel ndcontact -1322 467 -1322 467 1 nand21
rlabel pdcontact -1322 525 -1322 525 1 nand21
rlabel pdcontact -1351 524 -1351 524 1 nand21
rlabel polycontact -1300 484 -1300 484 1 nand21
rlabel polycontact -1304 590 -1304 590 1 nand22
rlabel ndcontact -1330 579 -1330 579 1 nand22
rlabel pdcontact -1347 626 -1347 626 1 nand22
rlabel polycontact -1354 598 -1354 598 1 p3
rlabel polycontact -1340 590 -1340 590 1 g2
rlabel metal1 -1290 590 -1290 590 1 p3g2
rlabel pdcontact -1297 609 -1297 609 1 p3g2
rlabel ndcontact -1297 582 -1297 582 1 p3g2
rlabel polycontact -1361 497 -1361 497 1 p3
rlabel polycontact -1348 489 -1348 489 1 p2
rlabel polycontact -1332 481 -1332 481 1 g1
rlabel metal1 -1286 484 -1286 484 1 p3p2g1
rlabel ndcontact -1293 476 -1293 476 1 p3p2g1
rlabel pdcontact -1293 503 -1293 503 1 p3p2g1
rlabel polycontact -1364 375 -1364 375 1 p3
rlabel polycontact -1351 367 -1351 367 1 p2
rlabel polycontact -1339 361 -1339 361 1 p1
rlabel polycontact -1328 356 -1328 356 1 g0
rlabel metal1 -1289 362 -1289 362 1 p3p2p1g0
rlabel ndcontact -1296 354 -1296 354 1 p3p2p1g0
rlabel pdcontact -1296 381 -1296 381 1 p3p2p1g0
rlabel polycontact -1231 498 -1231 498 1 p3g2
rlabel polycontact -1220 491 -1220 491 1 p3p2g1
rlabel polycontact -1209 484 -1209 484 1 p3p2p1g0
rlabel polycontact -1199 485 -1199 485 1 g3
rlabel metal1 -1007 43 -1007 43 5 vdd
rlabel pdcontact -1011 30 -1011 30 1 vdd
rlabel ndcontact -1011 3 -1011 3 1 gnd
rlabel metal1 -1009 -10 -1009 -10 1 gnd
rlabel metal1 -974 44 -974 44 5 vdd
rlabel pdcontact -978 31 -978 31 1 vdd
rlabel ndcontact -978 4 -978 4 1 gnd
rlabel metal1 -976 -9 -976 -9 1 gnd
rlabel pdcontact -919 31 -919 31 1 vdd
rlabel pdcontact -950 32 -950 32 1 vdd
rlabel ndcontact -950 -12 -950 -12 1 gnd
rlabel metal1 -936 47 -936 47 5 vdd
rlabel metal1 -892 -25 -892 -25 1 gnd
rlabel ndcontact -894 -12 -894 -12 1 gnd
rlabel pdcontact -894 15 -894 15 1 vdd
rlabel pdcontact -833 31 -833 31 1 vdd
rlabel pdcontact -864 32 -864 32 1 vdd
rlabel ndcontact -864 -12 -864 -12 1 gnd
rlabel metal1 -850 47 -850 47 5 vdd
rlabel metal1 -806 -25 -806 -25 1 gnd
rlabel ndcontact -808 -12 -808 -12 1 gnd
rlabel pdcontact -808 15 -808 15 1 vdd
rlabel pdcontact -740 17 -740 17 1 vdd
rlabel ndcontact -740 -10 -740 -10 1 gnd
rlabel metal1 -769 -27 -769 -27 1 gnd
rlabel metal1 -769 38 -769 38 5 vdd
rlabel pdcontact -778 20 -778 20 1 vdd
rlabel ndcontact -760 -17 -760 -17 1 gnd
rlabel ndcontact -778 -16 -778 -16 1 gnd
rlabel metal1 -1007 160 -1007 160 5 vdd
rlabel pdcontact -1011 147 -1011 147 1 vdd
rlabel ndcontact -1011 120 -1011 120 1 gnd
rlabel metal1 -1009 107 -1009 107 1 gnd
rlabel metal1 -974 161 -974 161 5 vdd
rlabel pdcontact -978 148 -978 148 1 vdd
rlabel ndcontact -978 121 -978 121 1 gnd
rlabel metal1 -976 108 -976 108 1 gnd
rlabel pdcontact -919 148 -919 148 1 vdd
rlabel pdcontact -950 149 -950 149 1 vdd
rlabel ndcontact -950 105 -950 105 1 gnd
rlabel metal1 -936 164 -936 164 5 vdd
rlabel metal1 -892 92 -892 92 1 gnd
rlabel ndcontact -894 105 -894 105 1 gnd
rlabel pdcontact -894 132 -894 132 1 vdd
rlabel pdcontact -833 148 -833 148 1 vdd
rlabel pdcontact -864 149 -864 149 1 vdd
rlabel ndcontact -864 105 -864 105 1 gnd
rlabel metal1 -850 164 -850 164 5 vdd
rlabel metal1 -806 92 -806 92 1 gnd
rlabel ndcontact -808 105 -808 105 1 gnd
rlabel pdcontact -808 132 -808 132 1 vdd
rlabel pdcontact -740 134 -740 134 1 vdd
rlabel ndcontact -740 107 -740 107 1 gnd
rlabel metal1 -769 90 -769 90 1 gnd
rlabel metal1 -769 155 -769 155 5 vdd
rlabel pdcontact -778 137 -778 137 1 vdd
rlabel ndcontact -760 100 -760 100 1 gnd
rlabel ndcontact -778 101 -778 101 1 gnd
rlabel polycontact -1010 11 -1010 11 1 p0
rlabel metal1 -996 11 -996 11 1 p01
rlabel pdcontact -1003 30 -1003 30 1 p01
rlabel ndcontact -1003 3 -1003 3 1 p01
rlabel polycontact -977 12 -977 12 1 c0
rlabel metal1 -963 12 -963 12 1 c01
rlabel pdcontact -970 31 -970 31 1 c01
rlabel ndcontact -970 4 -970 4 1 c01
rlabel polycontact -943 4 -943 4 1 p0
rlabel polycontact -929 -4 -929 -4 1 c01
rlabel pdcontact -936 32 -936 32 1 nand9
rlabel ndcontact -919 -15 -919 -15 1 nand9
rlabel polycontact -893 -4 -893 -4 1 nand9
rlabel ndcontact -886 -12 -886 -12 1 p0c01
rlabel metal1 -879 -4 -879 -4 1 p0c01
rlabel pdcontact -886 15 -886 15 1 p0c01
rlabel polycontact -857 4 -857 4 1 p01
rlabel polycontact -843 -4 -843 -4 1 c0
rlabel pdcontact -850 32 -850 32 1 nand10
rlabel ndcontact -833 -15 -833 -15 1 nand10
rlabel polycontact -807 -4 -807 -4 1 nand10
rlabel pdcontact -800 15 -800 15 1 p01c0
rlabel ndcontact -800 -12 -800 -12 1 p01c0
rlabel metal1 -793 -4 -793 -4 1 p01c0
rlabel polycontact -777 -1 -777 -1 1 p0c01
rlabel polycontact -766 -1 -766 -1 1 p01c0
rlabel pdcontact -759 20 -759 20 1 nor5
rlabel ndcontact -769 -17 -769 -17 1 nor5
rlabel polycontact -739 -2 -739 -2 1 nor5
rlabel pdcontact -732 17 -732 17 1 s0
rlabel metal1 -725 -2 -725 -2 1 s0
rlabel ndcontact -732 -10 -732 -10 1 s0
rlabel ndiffusion -936 -15 -936 -15 1 n17
rlabel ndiffusion -850 -16 -850 -16 1 n18
rlabel pdiffusion -769 21 -769 21 1 n19
rlabel metal1 -725 115 -725 115 1 s1
rlabel ndcontact -732 107 -732 107 1 s1
rlabel pdcontact -732 134 -732 134 1 s1
rlabel polycontact -739 115 -739 115 1 nor6
rlabel pdcontact -759 137 -759 137 1 nor6
rlabel ndcontact -769 100 -769 100 1 nor6
rlabel polycontact -1010 128 -1010 128 1 p1
rlabel metal1 -996 128 -996 128 1 p11
rlabel pdcontact -1003 147 -1003 147 1 p11
rlabel ndcontact -1003 120 -1003 120 1 p11
rlabel metal1 -963 129 -963 129 1 c11
rlabel ndcontact -970 121 -970 121 1 c11
rlabel pdcontact -970 148 -970 148 1 c11
rlabel pdcontact -936 149 -936 149 1 nand11
rlabel ndcontact -919 102 -919 102 1 nand11
rlabel polycontact -893 113 -893 113 1 nand11
rlabel ndiffusion -936 102 -936 102 1 n20
rlabel ndiffusion -850 101 -850 101 1 n21
rlabel pdiffusion -769 138 -769 138 1 n22
rlabel polycontact -766 116 -766 116 1 p11c1
rlabel polycontact -777 116 -777 116 1 p1c11
rlabel metal1 -793 113 -793 113 1 p11c1
rlabel pdcontact -800 132 -800 132 1 p11c1
rlabel ndcontact -800 105 -800 105 1 p11c1
rlabel polycontact -807 113 -807 113 1 nand12
rlabel pdcontact -850 149 -850 149 1 nand12
rlabel ndcontact -833 102 -833 102 1 nand12
rlabel polycontact -857 121 -857 121 1 p11
rlabel ndcontact -886 105 -886 105 1 p1c11
rlabel metal1 -879 113 -879 113 1 p1c11
rlabel pdcontact -886 132 -886 132 1 p1c11
rlabel polycontact -929 113 -929 113 1 c11
rlabel polycontact -943 121 -943 121 1 p1
rlabel metal1 -1005 280 -1005 280 5 vdd
rlabel pdcontact -1009 267 -1009 267 1 vdd
rlabel ndcontact -1009 240 -1009 240 1 gnd
rlabel metal1 -1007 227 -1007 227 1 gnd
rlabel metal1 -972 281 -972 281 5 vdd
rlabel pdcontact -976 268 -976 268 1 vdd
rlabel ndcontact -976 241 -976 241 1 gnd
rlabel metal1 -974 228 -974 228 1 gnd
rlabel pdcontact -917 268 -917 268 1 vdd
rlabel pdcontact -948 269 -948 269 1 vdd
rlabel ndcontact -948 225 -948 225 1 gnd
rlabel metal1 -934 284 -934 284 5 vdd
rlabel metal1 -890 212 -890 212 1 gnd
rlabel ndcontact -892 225 -892 225 1 gnd
rlabel pdcontact -892 252 -892 252 1 vdd
rlabel pdcontact -831 268 -831 268 1 vdd
rlabel pdcontact -862 269 -862 269 1 vdd
rlabel ndcontact -862 225 -862 225 1 gnd
rlabel metal1 -848 284 -848 284 5 vdd
rlabel metal1 -804 212 -804 212 1 gnd
rlabel ndcontact -806 225 -806 225 1 gnd
rlabel pdcontact -806 252 -806 252 1 vdd
rlabel pdcontact -738 254 -738 254 1 vdd
rlabel ndcontact -738 227 -738 227 1 gnd
rlabel metal1 -767 210 -767 210 1 gnd
rlabel metal1 -767 275 -767 275 5 vdd
rlabel pdcontact -776 257 -776 257 1 vdd
rlabel ndcontact -758 220 -758 220 1 gnd
rlabel ndcontact -776 221 -776 221 1 gnd
rlabel metal1 -1005 397 -1005 397 5 vdd
rlabel pdcontact -1009 384 -1009 384 1 vdd
rlabel ndcontact -1009 357 -1009 357 1 gnd
rlabel metal1 -1007 344 -1007 344 1 gnd
rlabel metal1 -972 398 -972 398 5 vdd
rlabel pdcontact -976 385 -976 385 1 vdd
rlabel ndcontact -976 358 -976 358 1 gnd
rlabel metal1 -974 345 -974 345 1 gnd
rlabel pdcontact -917 385 -917 385 1 vdd
rlabel pdcontact -948 386 -948 386 1 vdd
rlabel ndcontact -948 342 -948 342 1 gnd
rlabel metal1 -934 401 -934 401 5 vdd
rlabel metal1 -890 329 -890 329 1 gnd
rlabel ndcontact -892 342 -892 342 1 gnd
rlabel pdcontact -892 369 -892 369 1 vdd
rlabel pdcontact -831 385 -831 385 1 vdd
rlabel pdcontact -862 386 -862 386 1 vdd
rlabel ndcontact -862 342 -862 342 1 gnd
rlabel metal1 -848 401 -848 401 5 vdd
rlabel metal1 -804 329 -804 329 1 gnd
rlabel ndcontact -806 342 -806 342 1 gnd
rlabel pdcontact -806 369 -806 369 1 vdd
rlabel pdcontact -738 371 -738 371 1 vdd
rlabel ndcontact -738 344 -738 344 1 gnd
rlabel metal1 -767 327 -767 327 1 gnd
rlabel metal1 -767 392 -767 392 5 vdd
rlabel pdcontact -776 374 -776 374 1 vdd
rlabel ndcontact -758 337 -758 337 1 gnd
rlabel ndcontact -776 338 -776 338 1 gnd
rlabel metal1 -723 235 -723 235 7 s2
rlabel ndcontact -730 227 -730 227 1 s2
rlabel pdcontact -730 254 -730 254 1 s2
rlabel polycontact -737 235 -737 235 1 nor7
rlabel pdcontact -757 257 -757 257 1 nor7
rlabel ndcontact -767 220 -767 220 1 nor7
rlabel polycontact -764 236 -764 236 1 p21c2
rlabel polycontact -775 236 -775 236 1 p2c21
rlabel ndiffusion -934 222 -934 222 1 n23
rlabel ndiffusion -848 221 -848 221 1 n24
rlabel pdiffusion -767 258 -767 258 1 n25
rlabel metal1 -791 233 -791 233 1 p21c2
rlabel pdcontact -934 269 -934 269 1 nand13
rlabel ndcontact -917 222 -917 222 1 nand13
rlabel polycontact -891 233 -891 233 1 nand13
rlabel polycontact -805 233 -805 233 1 nand14
rlabel ndcontact -831 222 -831 222 1 nand14
rlabel pdcontact -848 269 -848 269 1 nand14
rlabel ndcontact -798 225 -798 225 1 p21c2
rlabel pdcontact -798 252 -798 252 1 p21c2
rlabel polycontact -841 233 -841 233 1 c2
rlabel polycontact -855 241 -855 241 1 p21
rlabel metal1 -877 233 -877 233 1 p2c21
rlabel pdcontact -884 252 -884 252 1 p2c21
rlabel ndcontact -884 225 -884 225 1 p2c21
rlabel polycontact -927 233 -927 233 1 c21
rlabel polycontact -941 241 -941 241 1 p2
rlabel ndcontact -968 241 -968 241 1 c21
rlabel metal1 -961 249 -961 249 1 c21
rlabel pdcontact -968 268 -968 268 1 c21
rlabel polycontact -975 249 -975 249 1 c2
rlabel metal1 -994 248 -994 248 1 p21
rlabel polycontact -1008 248 -1008 248 1 p2
rlabel pdcontact -1001 267 -1001 267 1 p21
rlabel ndcontact -1001 240 -1001 240 1 p21
rlabel polycontact -737 352 -737 352 1 nor8
rlabel ndcontact -767 337 -767 337 1 nor8
rlabel pdcontact -757 374 -757 374 1 nor8
rlabel pdiffusion -767 375 -767 375 1 n26
rlabel ndiffusion -848 338 -848 338 1 n27
rlabel ndiffusion -934 339 -934 339 1 n28
rlabel ndcontact -917 339 -917 339 1 nand15
rlabel polycontact -891 350 -891 350 1 nand15
rlabel pdcontact -934 386 -934 386 1 nand15
rlabel ndcontact -831 339 -831 339 1 nand16
rlabel polycontact -805 350 -805 350 1 nand16
rlabel pdcontact -848 386 -848 386 1 nand16
rlabel metal1 -723 352 -723 352 7 s3
rlabel ndcontact -730 344 -730 344 1 s3
rlabel pdcontact -730 371 -730 371 1 s3
rlabel polycontact -1008 365 -1008 365 1 p3
rlabel metal1 -994 365 -994 365 1 p31
rlabel polycontact -975 366 -975 366 1 c3
rlabel ndcontact -1001 357 -1001 357 1 p31
rlabel pdcontact -1001 384 -1001 384 1 p31
rlabel metal1 -961 366 -961 366 1 c31
rlabel ndcontact -968 358 -968 358 1 c31
rlabel pdcontact -968 385 -968 385 1 c31
rlabel polycontact -941 358 -941 358 1 p3
rlabel polycontact -927 350 -927 350 1 c31
rlabel metal1 -877 350 -877 350 1 p3c31
rlabel ndcontact -884 342 -884 342 1 p3c31
rlabel pdcontact -884 369 -884 369 1 p3c31
rlabel polycontact -855 358 -855 358 1 p31
rlabel polycontact -841 350 -841 350 1 c3
rlabel metal1 -791 350 -791 350 1 p31c3
rlabel ndcontact -798 342 -798 342 1 p31c3
rlabel pdcontact -798 369 -798 369 1 p31c3
rlabel polycontact -775 353 -775 353 1 p3c31
rlabel polycontact -764 353 -764 353 1 p31c3
rlabel polycontact -977 129 -977 129 1 g0
rlabel polycontact -843 113 -843 113 1 g0
rlabel pdcontact -1648 24 -1648 24 1 vdd
rlabel ndcontact -1648 -3 -1648 -3 1 gnd
rlabel metal1 -1646 -16 -1646 -16 1 gnd
rlabel metal1 -1690 56 -1690 56 5 vdd
rlabel ndcontact -1704 -3 -1704 -3 1 gnd
rlabel pdcontact -1704 41 -1704 41 1 vdd
rlabel pdcontact -1673 40 -1673 40 1 vdd
rlabel polycontact -1697 13 -1697 13 1 a0
rlabel polycontact -1683 5 -1683 5 1 b0
rlabel pdcontact -1690 41 -1690 41 1 a0b0
rlabel ndcontact -1673 -6 -1673 -6 1 a0b0
rlabel polycontact -1647 5 -1647 5 1 a0b0
rlabel ndcontact -1640 -3 -1640 -3 1 g0
rlabel metal1 -1633 5 -1633 5 7 g0
rlabel pdcontact -1640 24 -1640 24 1 g0
rlabel metal1 -1893 140 -1893 140 5 vdd
rlabel pdcontact -1897 127 -1897 127 1 vdd
rlabel ndcontact -1897 100 -1897 100 1 gnd
rlabel metal1 -1895 87 -1895 87 1 gnd
rlabel metal1 -1860 141 -1860 141 5 vdd
rlabel pdcontact -1864 128 -1864 128 1 vdd
rlabel ndcontact -1864 101 -1864 101 1 gnd
rlabel metal1 -1862 88 -1862 88 1 gnd
rlabel ndiffusion -1822 82 -1822 82 1 n1
rlabel pdcontact -1805 128 -1805 128 1 vdd
rlabel pdcontact -1836 129 -1836 129 1 vdd
rlabel ndcontact -1836 85 -1836 85 1 gnd
rlabel metal1 -1822 144 -1822 144 5 vdd
rlabel metal1 -1778 72 -1778 72 1 gnd
rlabel ndcontact -1780 85 -1780 85 1 gnd
rlabel pdcontact -1780 112 -1780 112 1 vdd
rlabel pdcontact -1719 128 -1719 128 1 vdd
rlabel pdcontact -1750 129 -1750 129 1 vdd
rlabel ndcontact -1750 85 -1750 85 1 gnd
rlabel metal1 -1736 144 -1736 144 5 vdd
rlabel metal1 -1692 72 -1692 72 1 gnd
rlabel ndcontact -1694 85 -1694 85 1 gnd
rlabel pdcontact -1694 112 -1694 112 1 vdd
rlabel polycontact -1779 93 -1779 93 1 nand1
rlabel pdcontact -1822 129 -1822 129 1 nand1
rlabel ndiffusion -1736 81 -1736 81 1 n2
rlabel ndcontact -1805 82 -1805 82 1 nand1
rlabel ndcontact -1719 82 -1719 82 1 nand2
rlabel pdcontact -1736 129 -1736 129 1 nand2
rlabel polycontact -1693 93 -1693 93 1 nand2
rlabel pdcontact -1626 114 -1626 114 1 vdd
rlabel ndcontact -1626 87 -1626 87 1 gnd
rlabel metal1 -1655 70 -1655 70 1 gnd
rlabel metal1 -1655 135 -1655 135 5 vdd
rlabel pdcontact -1664 117 -1664 117 1 vdd
rlabel ndcontact -1646 80 -1646 80 1 gnd
rlabel ndcontact -1664 81 -1664 81 1 gnd
rlabel pdiffusion -1655 118 -1655 118 1 n3
rlabel pdcontact -1645 117 -1645 117 1 nor
rlabel ndcontact -1655 80 -1655 80 1 nor
rlabel polycontact -1625 95 -1625 95 1 nor
rlabel polycontact -1896 108 -1896 108 1 a0
rlabel pdcontact -1889 127 -1889 127 1 a01
rlabel metal1 -1882 108 -1882 108 1 a01
rlabel ndcontact -1889 100 -1889 100 1 a01
rlabel polycontact -1863 109 -1863 109 1 b0
rlabel ndcontact -1856 101 -1856 101 1 b01
rlabel metal1 -1849 109 -1849 109 1 b01
rlabel pdcontact -1856 128 -1856 128 1 b01
rlabel polycontact -1829 101 -1829 101 1 a0
rlabel polycontact -1815 93 -1815 93 1 b01
rlabel pdcontact -1772 112 -1772 112 1 a0b01
rlabel metal1 -1765 93 -1765 93 1 a0b01
rlabel ndcontact -1772 85 -1772 85 1 a0b01
rlabel polycontact -1743 101 -1743 101 1 a01
rlabel polycontact -1729 93 -1729 93 1 b0
rlabel pdcontact -1686 112 -1686 112 1 a01b0
rlabel metal1 -1679 93 -1679 93 1 a01b0
rlabel ndcontact -1686 85 -1686 85 1 a01b0
rlabel polycontact -1663 96 -1663 96 1 a0b01
rlabel polycontact -1652 96 -1652 96 1 a01b0
rlabel ndiffusion -1690 -6 -1690 -6 1 n4
rlabel ndcontact -1618 87 -1618 87 1 p0
rlabel metal1 -1611 95 -1611 95 7 p0
rlabel pdcontact -1618 114 -1618 114 1 p0
rlabel pdcontact -1651 252 -1651 252 1 vdd
rlabel ndcontact -1651 225 -1651 225 1 gnd
rlabel metal1 -1649 212 -1649 212 1 gnd
rlabel metal1 -1693 284 -1693 284 5 vdd
rlabel ndcontact -1707 225 -1707 225 1 gnd
rlabel pdcontact -1707 269 -1707 269 1 vdd
rlabel pdcontact -1676 268 -1676 268 1 vdd
rlabel metal1 -1896 368 -1896 368 5 vdd
rlabel pdcontact -1900 355 -1900 355 1 vdd
rlabel ndcontact -1900 328 -1900 328 1 gnd
rlabel metal1 -1898 315 -1898 315 1 gnd
rlabel metal1 -1863 369 -1863 369 5 vdd
rlabel pdcontact -1867 356 -1867 356 1 vdd
rlabel ndcontact -1867 329 -1867 329 1 gnd
rlabel metal1 -1865 316 -1865 316 1 gnd
rlabel pdcontact -1808 356 -1808 356 1 vdd
rlabel pdcontact -1839 357 -1839 357 1 vdd
rlabel ndcontact -1839 313 -1839 313 1 gnd
rlabel metal1 -1825 372 -1825 372 5 vdd
rlabel metal1 -1781 300 -1781 300 1 gnd
rlabel ndcontact -1783 313 -1783 313 1 gnd
rlabel pdcontact -1783 340 -1783 340 1 vdd
rlabel pdcontact -1722 356 -1722 356 1 vdd
rlabel pdcontact -1753 357 -1753 357 1 vdd
rlabel ndcontact -1753 313 -1753 313 1 gnd
rlabel metal1 -1739 372 -1739 372 5 vdd
rlabel metal1 -1695 300 -1695 300 1 gnd
rlabel ndcontact -1697 313 -1697 313 1 gnd
rlabel pdcontact -1697 340 -1697 340 1 vdd
rlabel pdcontact -1629 342 -1629 342 1 vdd
rlabel ndcontact -1629 315 -1629 315 1 gnd
rlabel metal1 -1658 298 -1658 298 1 gnd
rlabel metal1 -1658 363 -1658 363 5 vdd
rlabel pdcontact -1667 345 -1667 345 1 vdd
rlabel ndcontact -1649 308 -1649 308 1 gnd
rlabel ndcontact -1667 309 -1667 309 1 gnd
rlabel pdcontact -1650 467 -1650 467 1 vdd
rlabel ndcontact -1650 440 -1650 440 1 gnd
rlabel metal1 -1648 427 -1648 427 1 gnd
rlabel metal1 -1692 499 -1692 499 5 vdd
rlabel ndcontact -1706 440 -1706 440 1 gnd
rlabel pdcontact -1706 484 -1706 484 1 vdd
rlabel pdcontact -1675 483 -1675 483 1 vdd
rlabel metal1 -1895 583 -1895 583 5 vdd
rlabel pdcontact -1899 570 -1899 570 1 vdd
rlabel ndcontact -1899 543 -1899 543 1 gnd
rlabel metal1 -1897 530 -1897 530 1 gnd
rlabel metal1 -1862 584 -1862 584 5 vdd
rlabel pdcontact -1866 571 -1866 571 1 vdd
rlabel ndcontact -1866 544 -1866 544 1 gnd
rlabel metal1 -1864 531 -1864 531 1 gnd
rlabel pdcontact -1807 571 -1807 571 1 vdd
rlabel pdcontact -1838 572 -1838 572 1 vdd
rlabel ndcontact -1838 528 -1838 528 1 gnd
rlabel metal1 -1824 587 -1824 587 5 vdd
rlabel metal1 -1780 515 -1780 515 1 gnd
rlabel ndcontact -1782 528 -1782 528 1 gnd
rlabel pdcontact -1782 555 -1782 555 1 vdd
rlabel pdcontact -1721 571 -1721 571 1 vdd
rlabel pdcontact -1752 572 -1752 572 1 vdd
rlabel ndcontact -1752 528 -1752 528 1 gnd
rlabel metal1 -1738 587 -1738 587 5 vdd
rlabel metal1 -1694 515 -1694 515 1 gnd
rlabel ndcontact -1696 528 -1696 528 1 gnd
rlabel pdcontact -1696 555 -1696 555 1 vdd
rlabel pdcontact -1628 557 -1628 557 1 vdd
rlabel ndcontact -1628 530 -1628 530 1 gnd
rlabel metal1 -1657 513 -1657 513 1 gnd
rlabel metal1 -1657 578 -1657 578 5 vdd
rlabel pdcontact -1666 560 -1666 560 1 vdd
rlabel ndcontact -1648 523 -1648 523 1 gnd
rlabel ndcontact -1666 524 -1666 524 1 gnd
rlabel pdcontact -1648 679 -1648 679 1 vdd
rlabel ndcontact -1648 652 -1648 652 1 gnd
rlabel metal1 -1646 639 -1646 639 1 gnd
rlabel metal1 -1690 711 -1690 711 5 vdd
rlabel ndcontact -1704 652 -1704 652 1 gnd
rlabel pdcontact -1704 696 -1704 696 1 vdd
rlabel pdcontact -1673 695 -1673 695 1 vdd
rlabel metal1 -1893 795 -1893 795 5 vdd
rlabel pdcontact -1897 782 -1897 782 1 vdd
rlabel ndcontact -1897 755 -1897 755 1 gnd
rlabel metal1 -1895 742 -1895 742 1 gnd
rlabel metal1 -1860 796 -1860 796 5 vdd
rlabel pdcontact -1864 783 -1864 783 1 vdd
rlabel ndcontact -1864 756 -1864 756 1 gnd
rlabel metal1 -1862 743 -1862 743 1 gnd
rlabel pdcontact -1805 783 -1805 783 1 vdd
rlabel pdcontact -1836 784 -1836 784 1 vdd
rlabel ndcontact -1836 740 -1836 740 1 gnd
rlabel metal1 -1822 799 -1822 799 5 vdd
rlabel metal1 -1778 727 -1778 727 1 gnd
rlabel ndcontact -1780 740 -1780 740 1 gnd
rlabel pdcontact -1780 767 -1780 767 1 vdd
rlabel pdcontact -1719 783 -1719 783 1 vdd
rlabel pdcontact -1750 784 -1750 784 1 vdd
rlabel ndcontact -1750 740 -1750 740 1 gnd
rlabel metal1 -1736 799 -1736 799 5 vdd
rlabel metal1 -1692 727 -1692 727 1 gnd
rlabel ndcontact -1694 740 -1694 740 1 gnd
rlabel pdcontact -1694 767 -1694 767 1 vdd
rlabel pdcontact -1626 769 -1626 769 1 vdd
rlabel ndcontact -1626 742 -1626 742 1 gnd
rlabel metal1 -1655 725 -1655 725 1 gnd
rlabel metal1 -1655 790 -1655 790 5 vdd
rlabel pdcontact -1664 772 -1664 772 1 vdd
rlabel ndcontact -1646 735 -1646 735 1 gnd
rlabel ndcontact -1664 736 -1664 736 1 gnd
rlabel polycontact -1700 241 -1700 241 1 a1
rlabel polycontact -1686 233 -1686 233 1 b1
rlabel pdcontact -1693 269 -1693 269 1 a1b1
rlabel ndcontact -1676 222 -1676 222 1 a1b1
rlabel polycontact -1650 233 -1650 233 1 a1b1
rlabel pdcontact -1643 252 -1643 252 1 g1
rlabel metal1 -1636 233 -1636 233 1 g1
rlabel ndcontact -1621 315 -1621 315 1 p1
rlabel metal1 -1614 323 -1614 323 1 p1
rlabel pdcontact -1621 342 -1621 342 1 p1
rlabel polycontact -1628 323 -1628 323 1 nor2
rlabel pdcontact -1648 345 -1648 345 1 nor2
rlabel ndcontact -1658 308 -1658 308 1 nor2
rlabel ndiffusion -1693 222 -1693 222 1 n5
rlabel pdiffusion -1658 346 -1658 346 1 n6
rlabel ndiffusion -1739 309 -1739 309 1 n7
rlabel ndiffusion -1825 310 -1825 310 1 n8
rlabel polycontact -1899 336 -1899 336 1 a1
rlabel metal1 -1885 336 -1885 336 1 a11
rlabel ndcontact -1892 328 -1892 328 1 a11
rlabel pdcontact -1892 355 -1892 355 1 a11
rlabel polycontact -1866 337 -1866 337 1 b1
rlabel metal1 -1852 337 -1852 337 1 b11
rlabel pdcontact -1859 356 -1859 356 1 b11
rlabel ndcontact -1859 329 -1859 329 1 b11
rlabel pdcontact -1825 357 -1825 357 1 nand3
rlabel ndcontact -1808 310 -1808 310 1 nand3
rlabel polycontact -1782 321 -1782 321 1 nand3
rlabel polycontact -1832 330 -1832 330 1 a1
rlabel polycontact -1818 321 -1818 321 1 b11
rlabel pdcontact -1775 340 -1775 340 1 a1b11
rlabel metal1 -1768 321 -1768 321 1 a1b11
rlabel ndcontact -1775 313 -1775 313 1 a1b11
rlabel polycontact -1746 329 -1746 329 1 a11
rlabel polycontact -1732 321 -1732 321 1 b1
rlabel pdcontact -1739 357 -1739 357 1 nand4
rlabel ndcontact -1722 310 -1722 310 1 nand4
rlabel polycontact -1696 321 -1696 321 1 nand4
rlabel ndcontact -1689 313 -1689 313 1 a11b1
rlabel metal1 -1682 321 -1682 321 1 a11b1
rlabel pdcontact -1689 340 -1689 340 1 a11b1
rlabel polycontact -1666 324 -1666 324 1 a1b11
rlabel polycontact -1655 324 -1655 324 1 a11b1
rlabel ndcontact -1642 440 -1642 440 1 g2
rlabel metal1 -1635 448 -1635 448 1 g2
rlabel pdcontact -1642 467 -1642 467 1 g2
rlabel polycontact -1649 448 -1649 448 1 a2b2
rlabel ndcontact -1675 437 -1675 437 1 a2b2
rlabel pdcontact -1692 484 -1692 484 1 a2b2
rlabel ndiffusion -1692 437 -1692 437 1 n9
rlabel polycontact -1685 448 -1685 448 1 b2
rlabel polycontact -1699 456 -1699 456 1 a2
rlabel polycontact -1627 538 -1627 538 1 nor3
rlabel pdiffusion -1657 561 -1657 561 1 n10
rlabel ndiffusion -1738 524 -1738 524 1 n11
rlabel ndiffusion -1824 525 -1824 525 1 n12
rlabel polycontact -1898 551 -1898 551 1 a2
rlabel metal1 -1884 551 -1884 551 1 a21
rlabel ndcontact -1891 543 -1891 543 1 a21
rlabel pdcontact -1891 570 -1891 570 1 a21
rlabel polycontact -1865 552 -1865 552 1 b2
rlabel pdcontact -1858 571 -1858 571 1 b21
rlabel metal1 -1851 552 -1851 552 1 b21
rlabel ndcontact -1858 544 -1858 544 1 b21
rlabel pdcontact -1824 572 -1824 572 1 nand5
rlabel polycontact -1831 544 -1831 544 1 a2
rlabel polycontact -1817 536 -1817 536 1 b21
rlabel ndcontact -1807 525 -1807 525 1 nand5
rlabel polycontact -1781 536 -1781 536 1 nand5
rlabel pdcontact -1774 555 -1774 555 1 a2b21
rlabel ndcontact -1774 528 -1774 528 1 a2b21
rlabel pdcontact -1738 572 -1738 572 1 nand6
rlabel ndcontact -1721 525 -1721 525 1 nand6
rlabel polycontact -1745 544 -1745 544 1 a21
rlabel polycontact -1731 536 -1731 536 1 b2
rlabel polycontact -1695 536 -1695 536 1 nand6
rlabel ndcontact -1688 528 -1688 528 1 a21b2
rlabel metal1 -1681 536 -1681 536 1 a21b2
rlabel pdcontact -1688 555 -1688 555 1 a21b2
rlabel metal1 -1767 536 -1767 536 1 a2b21
rlabel polycontact -1665 539 -1665 539 1 a2b21
rlabel polycontact -1654 539 -1654 539 1 a21b2
rlabel ndcontact -1657 523 -1657 523 1 nor3
rlabel pdcontact -1647 560 -1647 560 1 nor3
rlabel polycontact -1697 668 -1697 668 1 a3
rlabel polycontact -1683 660 -1683 660 1 b3
rlabel ndiffusion -1690 649 -1690 649 1 n13
rlabel pdcontact -1690 696 -1690 696 1 a3b3
rlabel ndcontact -1673 649 -1673 649 1 a3b3
rlabel polycontact -1647 660 -1647 660 1 a3b3
rlabel ndcontact -1640 652 -1640 652 1 g3
rlabel pdcontact -1640 679 -1640 679 1 g3
rlabel metal1 -1633 660 -1633 660 1 g3
rlabel metal1 -1611 750 -1611 750 7 p3
rlabel ndcontact -1618 742 -1618 742 1 p3
rlabel pdcontact -1618 769 -1618 769 1 p3
rlabel polycontact -1625 750 -1625 750 1 nor4
rlabel ndcontact -1655 735 -1655 735 1 nor4
rlabel pdcontact -1645 772 -1645 772 1 nor4
rlabel polycontact -1652 751 -1652 751 1 a31b3
rlabel polycontact -1663 751 -1663 751 1 a3b31
rlabel pdiffusion -1655 773 -1655 773 1 n14
rlabel ndcontact -1686 740 -1686 740 1 a31b3
rlabel metal1 -1679 748 -1679 748 1 a31b3
rlabel pdcontact -1686 767 -1686 767 1 a31b3
rlabel ndiffusion -1736 736 -1736 736 1 n15
rlabel ndiffusion -1822 737 -1822 737 1 n16
rlabel polycontact -1693 748 -1693 748 1 nand7
rlabel ndcontact -1719 737 -1719 737 1 nand7
rlabel pdcontact -1736 784 -1736 784 1 nand7
rlabel polycontact -1779 748 -1779 748 1 nand8
rlabel ndcontact -1805 737 -1805 737 1 nand8
rlabel pdcontact -1822 784 -1822 784 1 nand8
rlabel polycontact -1729 748 -1729 748 1 b3
rlabel polycontact -1743 756 -1743 756 1 a31
rlabel metal1 -1765 748 -1765 748 1 a3b31
rlabel pdcontact -1772 767 -1772 767 1 a3b31
rlabel ndcontact -1772 740 -1772 740 1 a3b31
rlabel polycontact -1829 756 -1829 756 1 a3
rlabel polycontact -1815 748 -1815 748 1 b31
rlabel metal1 -1849 764 -1849 764 1 b31
rlabel polycontact -1863 764 -1863 764 1 b3
rlabel pdcontact -1856 783 -1856 783 1 b31
rlabel ndcontact -1856 756 -1856 756 1 b31
rlabel polycontact -1896 763 -1896 763 1 a3
rlabel metal1 -1882 763 -1882 763 1 a31
rlabel ndcontact -1889 755 -1889 755 1 a31
rlabel pdcontact -1889 782 -1889 782 1 a31
rlabel ndcontact -1643 225 -1643 225 1 g1
rlabel ndcontact -1620 530 -1620 530 1 p2
rlabel metal1 -1613 538 -1613 538 1 p2
rlabel pdcontact -1620 557 -1620 557 1 p2
rlabel pdcontact -2179 -36 -2179 -36 1 vdd
rlabel polycontact -2168 -60 -2168 -60 1 clk
rlabel ndcontact -2179 -68 -2179 -68 1 gnd
rlabel pdcontact -2147 -36 -2147 -36 1 vdd
rlabel ndcontact -2147 -70 -2147 -70 1 gnd
rlabel ndcontact -2111 -70 -2111 -70 1 gnd
rlabel polycontact -2098 -60 -2098 -60 1 clk
rlabel pdcontact -2111 -37 -2111 -37 1 vdd
rlabel polycontact -2146 -56 -2146 -56 1 clk
rlabel metal1 -2058 -22 -2058 -22 5 vdd
rlabel pdcontact -2062 -35 -2062 -35 1 vdd
rlabel ndcontact -2062 -62 -2062 -62 1 gnd
rlabel metal1 -2060 -75 -2060 -75 1 gnd
rlabel pdcontact -2175 110 -2175 110 1 vdd
rlabel polycontact -2164 86 -2164 86 1 clk
rlabel ndcontact -2175 78 -2175 78 1 gnd
rlabel pdcontact -2143 110 -2143 110 1 vdd
rlabel ndcontact -2143 76 -2143 76 1 gnd
rlabel ndcontact -2107 76 -2107 76 1 gnd
rlabel polycontact -2094 86 -2094 86 1 clk
rlabel pdcontact -2107 109 -2107 109 1 vdd
rlabel polycontact -2142 90 -2142 90 1 clk
rlabel metal1 -2054 124 -2054 124 5 vdd
rlabel pdcontact -2058 111 -2058 111 1 vdd
rlabel ndcontact -2058 84 -2058 84 1 gnd
rlabel metal1 -2056 71 -2056 71 1 gnd
rlabel pdcontact -2181 238 -2181 238 1 vdd
rlabel polycontact -2170 214 -2170 214 1 clk
rlabel ndcontact -2181 206 -2181 206 1 gnd
rlabel pdcontact -2149 238 -2149 238 1 vdd
rlabel ndcontact -2149 204 -2149 204 1 gnd
rlabel ndcontact -2113 204 -2113 204 1 gnd
rlabel polycontact -2100 214 -2100 214 1 clk
rlabel pdcontact -2113 237 -2113 237 1 vdd
rlabel polycontact -2148 218 -2148 218 1 clk
rlabel metal1 -2060 252 -2060 252 5 vdd
rlabel pdcontact -2064 239 -2064 239 1 vdd
rlabel ndcontact -2064 212 -2064 212 1 gnd
rlabel metal1 -2062 199 -2062 199 1 gnd
rlabel pdcontact -2175 347 -2175 347 1 vdd
rlabel polycontact -2164 323 -2164 323 1 clk
rlabel ndcontact -2175 315 -2175 315 1 gnd
rlabel pdcontact -2143 347 -2143 347 1 vdd
rlabel ndcontact -2143 313 -2143 313 1 gnd
rlabel ndcontact -2107 313 -2107 313 1 gnd
rlabel polycontact -2094 323 -2094 323 1 clk
rlabel pdcontact -2107 346 -2107 346 1 vdd
rlabel polycontact -2142 327 -2142 327 1 clk
rlabel metal1 -2054 361 -2054 361 5 vdd
rlabel pdcontact -2058 348 -2058 348 1 vdd
rlabel ndcontact -2058 321 -2058 321 1 gnd
rlabel metal1 -2056 308 -2056 308 1 gnd
rlabel pdcontact -2167 455 -2167 455 1 vdd
rlabel polycontact -2156 431 -2156 431 1 clk
rlabel ndcontact -2167 423 -2167 423 1 gnd
rlabel pdcontact -2135 455 -2135 455 1 vdd
rlabel ndcontact -2135 421 -2135 421 1 gnd
rlabel ndcontact -2099 421 -2099 421 1 gnd
rlabel polycontact -2086 431 -2086 431 1 clk
rlabel pdcontact -2099 454 -2099 454 1 vdd
rlabel polycontact -2134 435 -2134 435 1 clk
rlabel metal1 -2046 469 -2046 469 5 vdd
rlabel pdcontact -2050 456 -2050 456 1 vdd
rlabel ndcontact -2050 429 -2050 429 1 gnd
rlabel metal1 -2048 416 -2048 416 1 gnd
rlabel pdcontact -2167 594 -2167 594 1 vdd
rlabel polycontact -2156 570 -2156 570 1 clk
rlabel ndcontact -2167 562 -2167 562 1 gnd
rlabel pdcontact -2135 594 -2135 594 1 vdd
rlabel ndcontact -2135 560 -2135 560 1 gnd
rlabel ndcontact -2099 560 -2099 560 1 gnd
rlabel polycontact -2086 570 -2086 570 1 clk
rlabel pdcontact -2099 593 -2099 593 1 vdd
rlabel polycontact -2134 574 -2134 574 1 clk
rlabel metal1 -2046 608 -2046 608 5 vdd
rlabel pdcontact -2050 595 -2050 595 1 vdd
rlabel ndcontact -2050 568 -2050 568 1 gnd
rlabel metal1 -2048 555 -2048 555 1 gnd
rlabel pdcontact -2154 719 -2154 719 1 vdd
rlabel polycontact -2143 695 -2143 695 1 clk
rlabel ndcontact -2154 687 -2154 687 1 gnd
rlabel pdcontact -2122 719 -2122 719 1 vdd
rlabel ndcontact -2122 685 -2122 685 1 gnd
rlabel ndcontact -2086 685 -2086 685 1 gnd
rlabel polycontact -2073 695 -2073 695 1 clk
rlabel pdcontact -2086 718 -2086 718 1 vdd
rlabel polycontact -2121 699 -2121 699 1 clk
rlabel metal1 -2033 733 -2033 733 5 vdd
rlabel pdcontact -2037 720 -2037 720 1 vdd
rlabel ndcontact -2037 693 -2037 693 1 gnd
rlabel metal1 -2035 680 -2035 680 1 gnd
rlabel pdcontact -2156 820 -2156 820 1 vdd
rlabel polycontact -2145 796 -2145 796 1 clk
rlabel ndcontact -2156 788 -2156 788 1 gnd
rlabel pdcontact -2124 820 -2124 820 1 vdd
rlabel ndcontact -2124 786 -2124 786 1 gnd
rlabel ndcontact -2088 786 -2088 786 1 gnd
rlabel polycontact -2075 796 -2075 796 1 clk
rlabel pdcontact -2088 819 -2088 819 1 vdd
rlabel polycontact -2123 800 -2123 800 1 clk
rlabel metal1 -2035 834 -2035 834 5 vdd
rlabel pdcontact -2039 821 -2039 821 1 vdd
rlabel ndcontact -2039 794 -2039 794 1 gnd
rlabel metal1 -2037 781 -2037 781 1 gnd
rlabel pdcontact -2152 -164 -2152 -164 1 vdd
rlabel polycontact -2141 -188 -2141 -188 1 clk
rlabel ndcontact -2152 -196 -2152 -196 1 gnd
rlabel pdcontact -2120 -164 -2120 -164 1 vdd
rlabel ndcontact -2120 -198 -2120 -198 1 gnd
rlabel ndcontact -2084 -198 -2084 -198 1 gnd
rlabel polycontact -2071 -188 -2071 -188 1 clk
rlabel pdcontact -2084 -165 -2084 -165 1 vdd
rlabel polycontact -2119 -184 -2119 -184 1 clk
rlabel metal1 -2031 -150 -2031 -150 5 vdd
rlabel pdcontact -2035 -163 -2035 -163 1 vdd
rlabel ndcontact -2035 -190 -2035 -190 1 gnd
rlabel metal1 -2033 -203 -2033 -203 1 gnd
rlabel polycontact -2151 -184 -2151 -184 1 a_0
rlabel metal1 -2020 -182 -2020 -182 1 a0
rlabel ndcontact -2027 -190 -2027 -190 1 a0
rlabel pdcontact -2027 -163 -2027 -163 1 a0
rlabel pdiffusion -2144 -164 -2144 -164 1 n45
rlabel ndiffusion -2111 -198 -2111 -198 1 n46
rlabel ndiffusion -2074 -198 -2074 -198 1 n47
rlabel polycontact -2034 -182 -2034 -182 1 n48
rlabel pdcontact -2061 -164 -2061 -164 1 n48
rlabel ndcontact -2061 -198 -2061 -198 1 n48
rlabel pdcontact -2132 -164 -2132 -164 1 x1
rlabel ndcontact -2132 -196 -2132 -196 1 x1
rlabel polycontact -2108 -188 -2108 -188 1 x1
rlabel polycontact -2082 -184 -2082 -184 1 y1
rlabel ndcontact -2097 -198 -2097 -198 1 y1
rlabel pdcontact -2097 -164 -2097 -164 1 y1
rlabel polycontact -2178 -56 -2178 -56 1 b_0
rlabel ndcontact -2159 -68 -2159 -68 1 x2
rlabel polycontact -2135 -60 -2135 -60 1 x2
rlabel pdcontact -2159 -36 -2159 -36 1 x2
rlabel pdcontact -2124 -36 -2124 -36 1 y2
rlabel polycontact -2109 -56 -2109 -56 1 y2
rlabel ndcontact -2124 -70 -2124 -70 1 y2
rlabel ndcontact -2054 -62 -2054 -62 1 b0
rlabel metal1 -2047 -54 -2047 -54 1 b0
rlabel pdcontact -2054 -35 -2054 -35 1 b0
rlabel pdiffusion -2171 -36 -2171 -36 1 n49
rlabel ndiffusion -2138 -70 -2138 -70 1 n50
rlabel ndiffusion -2100 -70 -2100 -70 1 n51
rlabel ndcontact -2088 -70 -2088 -70 1 n52
rlabel pdcontact -2088 -36 -2088 -36 1 n52
rlabel polycontact -2061 -54 -2061 -54 1 n52
rlabel pdiffusion -2167 110 -2167 110 1 n53
rlabel ndiffusion -2134 76 -2134 76 1 n54
rlabel ndiffusion -2097 76 -2097 76 1 n55
rlabel ndcontact -2084 76 -2084 76 1 n56
rlabel pdcontact -2084 110 -2084 110 1 n56
rlabel polycontact -2057 92 -2057 92 1 n56
rlabel ndcontact -2050 84 -2050 84 1 a1
rlabel metal1 -2043 92 -2043 92 1 a1
rlabel pdcontact -2050 111 -2050 111 1 a1
rlabel polycontact -2174 90 -2174 90 1 a_1
rlabel ndcontact -2155 78 -2155 78 1 x3
rlabel polycontact -2131 86 -2131 86 1 x3
rlabel pdcontact -2155 110 -2155 110 1 x3
rlabel polycontact -2105 90 -2105 90 1 y3
rlabel pdcontact -2120 110 -2120 110 1 y3
rlabel ndcontact -2120 76 -2120 76 1 y3
rlabel pdiffusion -2173 238 -2173 238 1 n57
rlabel ndiffusion -2140 204 -2140 204 1 n58
rlabel ndiffusion -2103 204 -2103 204 1 n59
rlabel ndcontact -2090 204 -2090 204 1 n60
rlabel pdcontact -2090 238 -2090 238 1 n60
rlabel polycontact -2063 220 -2063 220 1 n60
rlabel metal1 -2049 220 -2049 220 1 b1
rlabel ndcontact -2056 212 -2056 212 1 b1
rlabel pdcontact -2056 239 -2056 239 1 b1
rlabel polycontact -2180 218 -2180 218 1 b_1
rlabel pdcontact -2161 238 -2161 238 1 x4
rlabel ndcontact -2161 206 -2161 206 1 x4
rlabel polycontact -2137 214 -2137 214 1 x4
rlabel pdcontact -2126 238 -2126 238 1 y4
rlabel polycontact -2111 218 -2111 218 1 y4
rlabel ndcontact -2126 204 -2126 204 1 y4
rlabel pdiffusion -2167 347 -2167 347 1 n61
rlabel ndiffusion -2134 313 -2134 313 1 n62
rlabel ndiffusion -2097 313 -2097 313 1 n63
rlabel ndcontact -2084 313 -2084 313 1 n64
rlabel pdcontact -2084 345 -2084 345 1 n64
rlabel polycontact -2057 329 -2057 329 1 n64
rlabel metal1 -2043 329 -2043 329 1 a2
rlabel ndcontact -2050 321 -2050 321 1 a2
rlabel pdcontact -2050 348 -2050 348 1 a2
rlabel polycontact -2105 327 -2105 327 1 y5
rlabel pdcontact -2120 347 -2120 347 1 y5
rlabel ndcontact -2120 313 -2120 313 1 y5
rlabel polycontact -2131 323 -2131 323 1 x5
rlabel pdcontact -2155 347 -2155 347 1 x5
rlabel ndcontact -2155 315 -2155 315 1 x5
rlabel polycontact -2174 327 -2174 327 1 a_2
rlabel polycontact -2166 435 -2166 435 1 b_2
rlabel pdiffusion -2159 455 -2159 455 1 n65
rlabel ndiffusion -2126 421 -2126 421 1 n66
rlabel ndiffusion -2089 421 -2089 421 1 n67
rlabel ndcontact -2076 421 -2076 421 1 n68
rlabel pdcontact -2076 455 -2076 455 1 n68
rlabel polycontact -2049 437 -2049 437 1 n68
rlabel pdcontact -2042 456 -2042 456 1 b2
rlabel metal1 -2035 437 -2035 437 1 b2
rlabel ndcontact -2042 429 -2042 429 1 b2
rlabel polycontact -2097 435 -2097 435 1 y6
rlabel ndcontact -2112 421 -2112 421 1 y6
rlabel pdcontact -2112 455 -2112 455 1 y6
rlabel polycontact -2123 431 -2123 431 1 x6
rlabel ndcontact -2147 423 -2147 423 1 x6
rlabel pdcontact -2147 455 -2147 455 1 x6
rlabel pdiffusion -2159 594 -2159 594 1 n69
rlabel ndiffusion -2126 560 -2126 560 1 n70
rlabel ndiffusion -2088 560 -2088 560 1 n71
rlabel ndcontact -2076 560 -2076 560 1 n72
rlabel pdcontact -2076 594 -2076 594 1 n72
rlabel polycontact -2049 576 -2049 576 1 n72
rlabel metal1 -2035 576 -2035 576 1 a3
rlabel ndcontact -2042 568 -2042 568 1 a3
rlabel pdcontact -2042 595 -2042 595 1 a3
rlabel polycontact -2097 574 -2097 574 1 y7
rlabel ndcontact -2112 560 -2112 560 1 y7
rlabel pdcontact -2112 594 -2112 594 1 y7
rlabel polycontact -2123 570 -2123 570 1 x7
rlabel polycontact -2166 574 -2166 574 1 a_3
rlabel pdiffusion -2146 719 -2146 719 1 n73
rlabel ndiffusion -2113 685 -2113 685 1 n74
rlabel ndiffusion -2076 685 -2076 685 1 n75
rlabel ndcontact -2063 685 -2063 685 1 n76
rlabel pdcontact -2063 719 -2063 719 1 n76
rlabel polycontact -2036 701 -2036 701 1 n76
rlabel metal1 -2022 701 -2022 701 1 b3
rlabel ndcontact -2029 693 -2029 693 1 b3
rlabel pdcontact -2029 720 -2029 720 1 b3
rlabel polycontact -2084 699 -2084 699 1 y8
rlabel ndcontact -2099 685 -2099 685 1 y8
rlabel pdcontact -2099 719 -2099 719 1 y8
rlabel polycontact -2110 695 -2110 695 1 x8
rlabel pdcontact -2134 719 -2134 719 1 x8
rlabel ndcontact -2134 687 -2134 687 1 x8
rlabel polycontact -2153 699 -2153 699 1 b_3
rlabel pdiffusion -2148 820 -2148 820 1 n77
rlabel ndiffusion -2115 786 -2115 786 1 n78
rlabel ndiffusion -2078 786 -2078 786 1 n79
rlabel ndcontact -2065 786 -2065 786 1 n80
rlabel pdcontact -2065 820 -2065 820 1 n80
rlabel polycontact -2038 802 -2038 802 1 n80
rlabel metal1 -2024 802 -2024 802 1 c0
rlabel ndcontact -2031 794 -2031 794 1 c0
rlabel pdcontact -2031 821 -2031 821 1 c0
rlabel polycontact -2086 800 -2086 800 1 y9
rlabel ndcontact -2101 786 -2101 786 1 y9
rlabel pdcontact -2101 820 -2101 820 1 y9
rlabel polycontact -2112 796 -2112 796 1 x9
rlabel ndcontact -2136 788 -2136 788 1 x9
rlabel pdcontact -2136 820 -2136 820 1 x9
rlabel polycontact -2155 800 -2155 800 1 cin
rlabel pdcontact -561 -1 -561 -1 1 vdd
rlabel polycontact -550 -25 -550 -25 1 clk
rlabel ndcontact -561 -33 -561 -33 1 gnd
rlabel pdcontact -529 -1 -529 -1 1 vdd
rlabel ndcontact -529 -35 -529 -35 1 gnd
rlabel ndcontact -493 -35 -493 -35 1 gnd
rlabel polycontact -480 -25 -480 -25 1 clk
rlabel pdcontact -493 -2 -493 -2 1 vdd
rlabel polycontact -528 -21 -528 -21 1 clk
rlabel metal1 -440 13 -440 13 5 vdd
rlabel pdcontact -444 0 -444 0 1 vdd
rlabel ndcontact -444 -27 -444 -27 1 gnd
rlabel metal1 -442 -40 -442 -40 1 gnd
rlabel pdcontact -553 107 -553 107 1 vdd
rlabel polycontact -542 83 -542 83 1 clk
rlabel ndcontact -553 75 -553 75 1 gnd
rlabel pdcontact -521 107 -521 107 1 vdd
rlabel ndcontact -521 73 -521 73 1 gnd
rlabel ndcontact -485 73 -485 73 1 gnd
rlabel polycontact -472 83 -472 83 1 clk
rlabel pdcontact -485 106 -485 106 1 vdd
rlabel polycontact -520 87 -520 87 1 clk
rlabel metal1 -432 121 -432 121 5 vdd
rlabel pdcontact -436 108 -436 108 1 vdd
rlabel ndcontact -436 81 -436 81 1 gnd
rlabel metal1 -434 68 -434 68 1 gnd
rlabel pdcontact -553 246 -553 246 1 vdd
rlabel polycontact -542 222 -542 222 1 clk
rlabel ndcontact -553 214 -553 214 1 gnd
rlabel pdcontact -521 246 -521 246 1 vdd
rlabel ndcontact -521 212 -521 212 1 gnd
rlabel ndcontact -485 212 -485 212 1 gnd
rlabel polycontact -472 222 -472 222 1 clk
rlabel pdcontact -485 245 -485 245 1 vdd
rlabel polycontact -520 226 -520 226 1 clk
rlabel metal1 -432 260 -432 260 5 vdd
rlabel pdcontact -436 247 -436 247 1 vdd
rlabel ndcontact -436 220 -436 220 1 gnd
rlabel metal1 -434 207 -434 207 1 gnd
rlabel pdcontact -540 371 -540 371 1 vdd
rlabel polycontact -529 347 -529 347 1 clk
rlabel ndcontact -540 339 -540 339 1 gnd
rlabel pdcontact -508 371 -508 371 1 vdd
rlabel ndcontact -508 337 -508 337 1 gnd
rlabel ndcontact -472 337 -472 337 1 gnd
rlabel polycontact -459 347 -459 347 1 clk
rlabel pdcontact -472 370 -472 370 1 vdd
rlabel polycontact -507 351 -507 351 1 clk
rlabel metal1 -419 385 -419 385 5 vdd
rlabel pdcontact -423 372 -423 372 1 vdd
rlabel ndcontact -423 345 -423 345 1 gnd
rlabel metal1 -421 332 -421 332 1 gnd
rlabel pdcontact -542 472 -542 472 1 vdd
rlabel polycontact -531 448 -531 448 1 clk
rlabel ndcontact -542 440 -542 440 1 gnd
rlabel pdcontact -510 472 -510 472 1 vdd
rlabel ndcontact -510 438 -510 438 1 gnd
rlabel ndcontact -474 438 -474 438 1 gnd
rlabel polycontact -461 448 -461 448 1 clk
rlabel pdcontact -474 471 -474 471 1 vdd
rlabel polycontact -509 452 -509 452 1 clk
rlabel metal1 -421 486 -421 486 5 vdd
rlabel pdcontact -425 473 -425 473 1 vdd
rlabel ndcontact -425 446 -425 446 1 gnd
rlabel metal1 -423 433 -423 433 1 gnd
rlabel polycontact -560 -21 -560 -21 1 s0
rlabel pdiffusion -553 -1 -553 -1 1 n81
rlabel ndiffusion -520 -35 -520 -35 1 n82
rlabel ndiffusion -483 -35 -483 -35 1 n83
rlabel ndcontact -470 -35 -470 -35 1 n84
rlabel pdcontact -470 -3 -470 -3 1 n84
rlabel polycontact -443 -19 -443 -19 1 n84
rlabel metal1 -429 -19 -429 -19 1 s_0
rlabel ndcontact -436 -27 -436 -27 1 s_0
rlabel pdcontact -436 0 -436 0 1 s_0
rlabel polycontact -491 -21 -491 -21 1 y10
rlabel pdcontact -506 -1 -506 -1 1 y10
rlabel ndcontact -506 -35 -506 -35 1 y10
rlabel polycontact -517 -25 -517 -25 1 x10
rlabel pdcontact -541 -1 -541 -1 1 x10
rlabel ndcontact -541 -33 -541 -33 1 x10
rlabel polycontact -552 87 -552 87 1 s1
rlabel pdiffusion -545 107 -545 107 1 n85
rlabel ndiffusion -512 73 -512 73 1 n86
rlabel ndiffusion -475 73 -475 73 1 n87
rlabel ndcontact -462 73 -462 73 1 n88
rlabel pdcontact -462 107 -462 107 1 n88
rlabel polycontact -435 89 -435 89 1 n88
rlabel ndcontact -428 81 -428 81 1 s_1
rlabel metal1 -421 89 -421 89 1 s_1
rlabel pdcontact -428 108 -428 108 1 s_1
rlabel polycontact -483 87 -483 87 1 y11
rlabel pdcontact -498 107 -498 107 1 y11
rlabel ndcontact -498 73 -498 73 1 y11
rlabel polycontact -509 83 -509 83 1 x11
rlabel pdcontact -533 107 -533 107 1 x11
rlabel ndcontact -533 75 -533 75 1 x11
rlabel polycontact -552 226 -552 226 1 s2
rlabel ndcontact -2147 562 -2147 562 1 x7
rlabel pdcontact -2147 594 -2147 594 1 x7
rlabel ndcontact -533 214 -533 214 1 x12
rlabel pdcontact -533 246 -533 246 1 x12
rlabel polycontact -509 222 -509 222 1 x12
rlabel pdiffusion -545 246 -545 246 1 n89
rlabel ndiffusion -512 212 -512 212 1 n90
rlabel ndiffusion -474 212 -474 212 1 n91
rlabel ndcontact -462 212 -462 212 1 n92
rlabel pdcontact -462 246 -462 246 1 n92
rlabel polycontact -435 228 -435 228 1 n92
rlabel polycontact -483 226 -483 226 1 y12
rlabel ndcontact -498 212 -498 212 1 y12
rlabel pdcontact -498 246 -498 246 1 y12
rlabel metal1 -421 228 -421 228 1 s_2
rlabel pdcontact -428 247 -428 247 1 s_2
rlabel ndcontact -428 220 -428 220 1 s_2
rlabel metal1 -408 353 -408 353 7 s_3
rlabel pdcontact -415 372 -415 372 1 s_3
rlabel ndcontact -415 345 -415 345 1 s_3
rlabel polycontact -422 353 -422 353 1 n96
rlabel ndcontact -449 337 -449 337 1 n96
rlabel pdcontact -449 371 -449 371 1 n96
rlabel ndiffusion -462 337 -462 337 1 n95
rlabel ndiffusion -499 337 -499 337 1 n94
rlabel pdiffusion -532 371 -532 371 1 n93
rlabel polycontact -539 351 -539 351 1 s3
rlabel ndcontact -520 339 -520 339 1 x13
rlabel pdcontact -520 371 -520 371 1 x13
rlabel polycontact -496 347 -496 347 1 x13
rlabel pdcontact -485 371 -485 371 1 y13
rlabel ndcontact -485 337 -485 337 1 y13
rlabel polycontact -470 351 -470 351 1 y13
rlabel polycontact -541 452 -541 452 1 c4
rlabel pdiffusion -534 472 -534 472 1 n97
rlabel ndiffusion -501 438 -501 438 1 n98
rlabel ndiffusion -464 438 -464 438 1 n99
rlabel ndcontact -451 438 -451 438 1 n100
rlabel pdcontact -451 472 -451 472 1 n100
rlabel polycontact -424 454 -424 454 1 n100
rlabel metal1 -410 454 -410 454 7 cout
rlabel ndcontact -417 446 -417 446 1 cout
rlabel pdcontact -417 473 -417 473 1 cout
rlabel polycontact -472 452 -472 452 1 y14
rlabel pdcontact -487 472 -487 472 1 y14
rlabel ndcontact -487 438 -487 438 1 y14
rlabel polycontact -498 448 -498 448 1 x14
rlabel pdcontact -522 472 -522 472 1 x14
rlabel ndcontact -522 440 -522 440 1 x14
<< end >>
